module font_rom(
input clk,
input [11:0] address,
output [7:0] out);

reg [7:0] font_rom [11:0];
reg [7:0] out;

//Source file: Untitled.raw
//Size: 65536 bytes

//Output file: Untitled.raw.dat
//ASCII 0x00 ' '
font_rom[0] <= 8'b00000000;
font_rom[1] <= 8'b00000000;
font_rom[2] <= 8'b00000000;
font_rom[3] <= 8'b00000000;
font_rom[4] <= 8'b00000000;
font_rom[5] <= 8'b00000000;
font_rom[6] <= 8'b00000000;
font_rom[7] <= 8'b00000000;
font_rom[8] <= 8'b00000000;
font_rom[9] <= 8'b00000000;
font_rom[10] <= 8'b00000000;
font_rom[11] <= 8'b00000000;
font_rom[12] <= 8'b00000000;
font_rom[13] <= 8'b00000000;
font_rom[14] <= 8'b00000000;
font_rom[15] <= 8'b00000000;
font_rom[16] <= 8'b00000000;
font_rom[17] <= 8'b00000000;
font_rom[18] <= 8'b00000000;
font_rom[19] <= 8'b00000000;
font_rom[20] <= 8'b00000000;
font_rom[21] <= 8'b00000000;
font_rom[22] <= 8'b00000000;
font_rom[23] <= 8'b00000000;
font_rom[24] <= 8'b00000000;
font_rom[25] <= 8'b00000000;
font_rom[26] <= 8'b00000000;
font_rom[27] <= 8'b00000000;
font_rom[28] <= 8'b00000000;
font_rom[29] <= 8'b00000000;
font_rom[30] <= 8'b00000000;
font_rom[31] <= 8'b00000000;
//ASCII 0x01 ' '
font_rom[32] <= 8'b00000000;
font_rom[33] <= 8'b00000000;
font_rom[34] <= 8'b00000000;
font_rom[35] <= 8'b00000000;
font_rom[36] <= 8'b00000000;
font_rom[37] <= 8'b00000000;
font_rom[38] <= 8'b00000000;
font_rom[39] <= 8'b00000000;
font_rom[40] <= 8'b00000000;
font_rom[41] <= 8'b00000000;
font_rom[42] <= 8'b00000000;
font_rom[43] <= 8'b00000000;
font_rom[44] <= 8'b00000000;
font_rom[45] <= 8'b00000000;
font_rom[46] <= 8'b00000000;
font_rom[47] <= 8'b00000000;
font_rom[48] <= 8'b00000000;
font_rom[49] <= 8'b00000000;
font_rom[50] <= 8'b00000000;
font_rom[51] <= 8'b00000000;
font_rom[52] <= 8'b00000000;
font_rom[53] <= 8'b00000000;
font_rom[54] <= 8'b00000000;
font_rom[55] <= 8'b00000000;
font_rom[56] <= 8'b00000000;
font_rom[57] <= 8'b00000000;
font_rom[58] <= 8'b00000000;
font_rom[59] <= 8'b00000000;
font_rom[60] <= 8'b00000000;
font_rom[61] <= 8'b00000000;
font_rom[62] <= 8'b00000000;
font_rom[63] <= 8'b00000000;
//ASCII 0x02 ' '
font_rom[64] <= 8'b00000000;
font_rom[65] <= 8'b00000000;
font_rom[66] <= 8'b00000000;
font_rom[67] <= 8'b00000000;
font_rom[68] <= 8'b00000000;
font_rom[69] <= 8'b00000000;
font_rom[70] <= 8'b00000000;
font_rom[71] <= 8'b00000000;
font_rom[72] <= 8'b00000000;
font_rom[73] <= 8'b00000000;
font_rom[74] <= 8'b00000000;
font_rom[75] <= 8'b00000000;
font_rom[76] <= 8'b00000000;
font_rom[77] <= 8'b00000000;
font_rom[78] <= 8'b00000000;
font_rom[79] <= 8'b00000000;
font_rom[80] <= 8'b00000000;
font_rom[81] <= 8'b00000000;
font_rom[82] <= 8'b00000000;
font_rom[83] <= 8'b00000000;
font_rom[84] <= 8'b00000111;
font_rom[85] <= 8'b10000000;
font_rom[86] <= 8'b00000000;
font_rom[87] <= 8'b10000000;
font_rom[88] <= 8'b00000000;
font_rom[89] <= 8'b10000000;
font_rom[90] <= 8'b00000000;
font_rom[91] <= 8'b10000000;
font_rom[92] <= 8'b00000000;
font_rom[93] <= 8'b10000000;
font_rom[94] <= 8'b00000000;
font_rom[95] <= 8'b10000000;
//ASCII 0x03 ' '
font_rom[96] <= 8'b00000000;
font_rom[97] <= 8'b00000000;
font_rom[98] <= 8'b00000000;
font_rom[99] <= 8'b00000000;
font_rom[100] <= 8'b00000000;
font_rom[101] <= 8'b00000000;
font_rom[102] <= 8'b00000000;
font_rom[103] <= 8'b00000000;
font_rom[104] <= 8'b00000000;
font_rom[105] <= 8'b10000000;
font_rom[106] <= 8'b00000000;
font_rom[107] <= 8'b10000000;
font_rom[108] <= 8'b00000000;
font_rom[109] <= 8'b10000000;
font_rom[110] <= 8'b00000000;
font_rom[111] <= 8'b10000000;
font_rom[112] <= 8'b00000000;
font_rom[113] <= 8'b10000000;
font_rom[114] <= 8'b00000000;
font_rom[115] <= 8'b10000000;
font_rom[116] <= 8'b00000000;
font_rom[117] <= 8'b11100000;
font_rom[118] <= 8'b00000000;
font_rom[119] <= 8'b00000000;
font_rom[120] <= 8'b00000000;
font_rom[121] <= 8'b00000000;
font_rom[122] <= 8'b00000000;
font_rom[123] <= 8'b00000000;
font_rom[124] <= 8'b00000000;
font_rom[125] <= 8'b00000000;
font_rom[126] <= 8'b00000000;
font_rom[127] <= 8'b00000000;
//ASCII 0x04 ' '
font_rom[128] <= 8'b00000000;
font_rom[129] <= 8'b00000000;
font_rom[130] <= 8'b00000000;
font_rom[131] <= 8'b00000000;
font_rom[132] <= 8'b00000000;
font_rom[133] <= 8'b00000000;
font_rom[134] <= 8'b00000000;
font_rom[135] <= 8'b00000000;
font_rom[136] <= 8'b00000000;
font_rom[137] <= 8'b10000000;
font_rom[138] <= 8'b00000000;
font_rom[139] <= 8'b10000000;
font_rom[140] <= 8'b00000000;
font_rom[141] <= 8'b10000000;
font_rom[142] <= 8'b00000000;
font_rom[143] <= 8'b10000000;
font_rom[144] <= 8'b00000000;
font_rom[145] <= 8'b10000000;
font_rom[146] <= 8'b00000000;
font_rom[147] <= 8'b10000000;
font_rom[148] <= 8'b00000111;
font_rom[149] <= 8'b10000000;
font_rom[150] <= 8'b00000000;
font_rom[151] <= 8'b00000000;
font_rom[152] <= 8'b00000000;
font_rom[153] <= 8'b00000000;
font_rom[154] <= 8'b00000000;
font_rom[155] <= 8'b00000000;
font_rom[156] <= 8'b00000000;
font_rom[157] <= 8'b00000000;
font_rom[158] <= 8'b00000000;
font_rom[159] <= 8'b00000000;
//ASCII 0x05 ' '
font_rom[160] <= 8'b00000000;
font_rom[161] <= 8'b00000000;
font_rom[162] <= 8'b00000000;
font_rom[163] <= 8'b00000000;
font_rom[164] <= 8'b00000000;
font_rom[165] <= 8'b00000000;
font_rom[166] <= 8'b00000000;
font_rom[167] <= 8'b00000000;
font_rom[168] <= 8'b00000000;
font_rom[169] <= 8'b10000000;
font_rom[170] <= 8'b00000000;
font_rom[171] <= 8'b10000000;
font_rom[172] <= 8'b00000000;
font_rom[173] <= 8'b10000000;
font_rom[174] <= 8'b00000000;
font_rom[175] <= 8'b10000000;
font_rom[176] <= 8'b00000000;
font_rom[177] <= 8'b10000000;
font_rom[178] <= 8'b00000000;
font_rom[179] <= 8'b10000000;
font_rom[180] <= 8'b00000000;
font_rom[181] <= 8'b10000000;
font_rom[182] <= 8'b00000000;
font_rom[183] <= 8'b10000000;
font_rom[184] <= 8'b00000000;
font_rom[185] <= 8'b10000000;
font_rom[186] <= 8'b00000000;
font_rom[187] <= 8'b10000000;
font_rom[188] <= 8'b00000000;
font_rom[189] <= 8'b10000000;
font_rom[190] <= 8'b00000000;
font_rom[191] <= 8'b10000000;
//ASCII 0x06 ' '
font_rom[192] <= 8'b00000000;
font_rom[193] <= 8'b00000000;
font_rom[194] <= 8'b00000000;
font_rom[195] <= 8'b00000000;
font_rom[196] <= 8'b00000000;
font_rom[197] <= 8'b00000000;
font_rom[198] <= 8'b00000000;
font_rom[199] <= 8'b00000000;
font_rom[200] <= 8'b00000000;
font_rom[201] <= 8'b00000000;
font_rom[202] <= 8'b00000000;
font_rom[203] <= 8'b00000000;
font_rom[204] <= 8'b00000000;
font_rom[205] <= 8'b00000000;
font_rom[206] <= 8'b00000000;
font_rom[207] <= 8'b00000000;
font_rom[208] <= 8'b00000000;
font_rom[209] <= 8'b00000000;
font_rom[210] <= 8'b00000000;
font_rom[211] <= 8'b00000000;
font_rom[212] <= 8'b00000111;
font_rom[213] <= 8'b11100000;
font_rom[214] <= 8'b00000000;
font_rom[215] <= 8'b00000000;
font_rom[216] <= 8'b00000000;
font_rom[217] <= 8'b00000000;
font_rom[218] <= 8'b00000000;
font_rom[219] <= 8'b00000000;
font_rom[220] <= 8'b00000000;
font_rom[221] <= 8'b00000000;
font_rom[222] <= 8'b00000000;
font_rom[223] <= 8'b00000000;
//ASCII 0x07 ' '
font_rom[224] <= 8'b00000000;
font_rom[225] <= 8'b00000000;
font_rom[226] <= 8'b00000000;
font_rom[227] <= 8'b00000000;
font_rom[228] <= 8'b00000000;
font_rom[229] <= 8'b00000000;
font_rom[230] <= 8'b00000000;
font_rom[231] <= 8'b00000000;
font_rom[232] <= 8'b00000000;
font_rom[233] <= 8'b00000000;
font_rom[234] <= 8'b00000000;
font_rom[235] <= 8'b00000000;
font_rom[236] <= 8'b00000000;
font_rom[237] <= 8'b00000000;
font_rom[238] <= 8'b00000001;
font_rom[239] <= 8'b10000000;
font_rom[240] <= 8'b00000011;
font_rom[241] <= 8'b11000000;
font_rom[242] <= 8'b00000011;
font_rom[243] <= 8'b11000000;
font_rom[244] <= 8'b00000011;
font_rom[245] <= 8'b11000000;
font_rom[246] <= 8'b00000001;
font_rom[247] <= 8'b10000000;
font_rom[248] <= 8'b00000000;
font_rom[249] <= 8'b00000000;
font_rom[250] <= 8'b00000000;
font_rom[251] <= 8'b00000000;
font_rom[252] <= 8'b00000000;
font_rom[253] <= 8'b00000000;
font_rom[254] <= 8'b00000000;
font_rom[255] <= 8'b00000000;
//ASCII 0x08 ' '
font_rom[256] <= 8'b00000000;
font_rom[257] <= 8'b00000000;
font_rom[258] <= 8'b00000000;
font_rom[259] <= 8'b00000000;
font_rom[260] <= 8'b00000000;
font_rom[261] <= 8'b00000000;
font_rom[262] <= 8'b00000000;
font_rom[263] <= 8'b00000000;
font_rom[264] <= 8'b00000111;
font_rom[265] <= 8'b11100000;
font_rom[266] <= 8'b00000111;
font_rom[267] <= 8'b11100000;
font_rom[268] <= 8'b00000111;
font_rom[269] <= 8'b11100000;
font_rom[270] <= 8'b00000110;
font_rom[271] <= 8'b01100000;
font_rom[272] <= 8'b00000100;
font_rom[273] <= 8'b00100000;
font_rom[274] <= 8'b00000100;
font_rom[275] <= 8'b00100000;
font_rom[276] <= 8'b00000100;
font_rom[277] <= 8'b00100000;
font_rom[278] <= 8'b00000110;
font_rom[279] <= 8'b01100000;
font_rom[280] <= 8'b00000111;
font_rom[281] <= 8'b11100000;
font_rom[282] <= 8'b00000111;
font_rom[283] <= 8'b11100000;
font_rom[284] <= 8'b00000111;
font_rom[285] <= 8'b11100000;
font_rom[286] <= 8'b00000111;
font_rom[287] <= 8'b11100000;
//ASCII 0x09 ' '
font_rom[288] <= 8'b00000000;
font_rom[289] <= 8'b00000000;
font_rom[290] <= 8'b00000000;
font_rom[291] <= 8'b00000000;
font_rom[292] <= 8'b00000000;
font_rom[293] <= 8'b00000000;
font_rom[294] <= 8'b00000000;
font_rom[295] <= 8'b00000000;
font_rom[296] <= 8'b00000000;
font_rom[297] <= 8'b00000000;
font_rom[298] <= 8'b00000000;
font_rom[299] <= 8'b00000000;
font_rom[300] <= 8'b00000000;
font_rom[301] <= 8'b00000000;
font_rom[302] <= 8'b00000000;
font_rom[303] <= 8'b00000000;
font_rom[304] <= 8'b00000000;
font_rom[305] <= 8'b00000000;
font_rom[306] <= 8'b00000000;
font_rom[307] <= 8'b00000000;
font_rom[308] <= 8'b00000000;
font_rom[309] <= 8'b00000000;
font_rom[310] <= 8'b00000000;
font_rom[311] <= 8'b00000000;
font_rom[312] <= 8'b00000000;
font_rom[313] <= 8'b00000000;
font_rom[314] <= 8'b00000000;
font_rom[315] <= 8'b00000000;
font_rom[316] <= 8'b00000000;
font_rom[317] <= 8'b00000000;
font_rom[318] <= 8'b00000000;
font_rom[319] <= 8'b00000000;
//ASCII 0x0A ' '
font_rom[320] <= 8'b00000000;
font_rom[321] <= 8'b00000000;
font_rom[322] <= 8'b00000000;
font_rom[323] <= 8'b00000000;
font_rom[324] <= 8'b00000000;
font_rom[325] <= 8'b00000000;
font_rom[326] <= 8'b00000000;
font_rom[327] <= 8'b00000000;
font_rom[328] <= 8'b00000000;
font_rom[329] <= 8'b00000000;
font_rom[330] <= 8'b00000000;
font_rom[331] <= 8'b00000000;
font_rom[332] <= 8'b00000000;
font_rom[333] <= 8'b00000000;
font_rom[334] <= 8'b00000000;
font_rom[335] <= 8'b00000000;
font_rom[336] <= 8'b00000000;
font_rom[337] <= 8'b00000000;
font_rom[338] <= 8'b00000000;
font_rom[339] <= 8'b00000000;
font_rom[340] <= 8'b00000000;
font_rom[341] <= 8'b00000000;
font_rom[342] <= 8'b00000000;
font_rom[343] <= 8'b00000000;
font_rom[344] <= 8'b00000000;
font_rom[345] <= 8'b00000000;
font_rom[346] <= 8'b00000000;
font_rom[347] <= 8'b00000000;
font_rom[348] <= 8'b00000000;
font_rom[349] <= 8'b00000000;
font_rom[350] <= 8'b00000000;
font_rom[351] <= 8'b00000000;
//ASCII 0x0B ' '
font_rom[352] <= 8'b00000000;
font_rom[353] <= 8'b00000000;
font_rom[354] <= 8'b00000000;
font_rom[355] <= 8'b00000000;
font_rom[356] <= 8'b00000000;
font_rom[357] <= 8'b00000000;
font_rom[358] <= 8'b00000000;
font_rom[359] <= 8'b00000000;
font_rom[360] <= 8'b00000000;
font_rom[361] <= 8'b00000000;
font_rom[362] <= 8'b00000000;
font_rom[363] <= 8'b11100000;
font_rom[364] <= 8'b00000000;
font_rom[365] <= 8'b01100000;
font_rom[366] <= 8'b00000000;
font_rom[367] <= 8'b01100000;
font_rom[368] <= 8'b00000000;
font_rom[369] <= 8'b10100000;
font_rom[370] <= 8'b00000000;
font_rom[371] <= 8'b10000000;
font_rom[372] <= 8'b00000001;
font_rom[373] <= 8'b10000000;
font_rom[374] <= 8'b00000010;
font_rom[375] <= 8'b01000000;
font_rom[376] <= 8'b00000010;
font_rom[377] <= 8'b01000000;
font_rom[378] <= 8'b00000001;
font_rom[379] <= 8'b10000000;
font_rom[380] <= 8'b00000000;
font_rom[381] <= 8'b00000000;
font_rom[382] <= 8'b00000000;
font_rom[383] <= 8'b00000000;
//ASCII 0x0C ' '
font_rom[384] <= 8'b00000000;
font_rom[385] <= 8'b00000000;
font_rom[386] <= 8'b00000000;
font_rom[387] <= 8'b00000000;
font_rom[388] <= 8'b00000000;
font_rom[389] <= 8'b00000000;
font_rom[390] <= 8'b00000000;
font_rom[391] <= 8'b00000000;
font_rom[392] <= 8'b00000000;
font_rom[393] <= 8'b00000000;
font_rom[394] <= 8'b00000001;
font_rom[395] <= 8'b11000000;
font_rom[396] <= 8'b00000010;
font_rom[397] <= 8'b00100000;
font_rom[398] <= 8'b00000010;
font_rom[399] <= 8'b00100000;
font_rom[400] <= 8'b00000001;
font_rom[401] <= 8'b11000000;
font_rom[402] <= 8'b00000000;
font_rom[403] <= 8'b10000000;
font_rom[404] <= 8'b00000011;
font_rom[405] <= 8'b11100000;
font_rom[406] <= 8'b00000000;
font_rom[407] <= 8'b10000000;
font_rom[408] <= 8'b00000000;
font_rom[409] <= 8'b10000000;
font_rom[410] <= 8'b00000000;
font_rom[411] <= 8'b10000000;
font_rom[412] <= 8'b00000000;
font_rom[413] <= 8'b00000000;
font_rom[414] <= 8'b00000000;
font_rom[415] <= 8'b00000000;
//ASCII 0x0D ' '
font_rom[416] <= 8'b00000000;
font_rom[417] <= 8'b00000000;
font_rom[418] <= 8'b00000000;
font_rom[419] <= 8'b00000000;
font_rom[420] <= 8'b00000000;
font_rom[421] <= 8'b00000000;
font_rom[422] <= 8'b00000000;
font_rom[423] <= 8'b00000000;
font_rom[424] <= 8'b00000000;
font_rom[425] <= 8'b00000000;
font_rom[426] <= 8'b00000000;
font_rom[427] <= 8'b00000000;
font_rom[428] <= 8'b00000000;
font_rom[429] <= 8'b00000000;
font_rom[430] <= 8'b00000000;
font_rom[431] <= 8'b00000000;
font_rom[432] <= 8'b00000000;
font_rom[433] <= 8'b00000000;
font_rom[434] <= 8'b00000000;
font_rom[435] <= 8'b00000000;
font_rom[436] <= 8'b00000000;
font_rom[437] <= 8'b00000000;
font_rom[438] <= 8'b00000000;
font_rom[439] <= 8'b00000000;
font_rom[440] <= 8'b00000000;
font_rom[441] <= 8'b00000000;
font_rom[442] <= 8'b00000000;
font_rom[443] <= 8'b00000000;
font_rom[444] <= 8'b00000000;
font_rom[445] <= 8'b00000000;
font_rom[446] <= 8'b00000000;
font_rom[447] <= 8'b00000000;
//ASCII 0x0E ' '
font_rom[448] <= 8'b00000000;
font_rom[449] <= 8'b00000000;
font_rom[450] <= 8'b00000000;
font_rom[451] <= 8'b00000000;
font_rom[452] <= 8'b00000000;
font_rom[453] <= 8'b00000000;
font_rom[454] <= 8'b00000000;
font_rom[455] <= 8'b00000000;
font_rom[456] <= 8'b00000000;
font_rom[457] <= 8'b00000000;
font_rom[458] <= 8'b00000000;
font_rom[459] <= 8'b01100000;
font_rom[460] <= 8'b00000001;
font_rom[461] <= 8'b10100000;
font_rom[462] <= 8'b00000001;
font_rom[463] <= 8'b01100000;
font_rom[464] <= 8'b00000001;
font_rom[465] <= 8'b10100000;
font_rom[466] <= 8'b00000001;
font_rom[467] <= 8'b00100000;
font_rom[468] <= 8'b00000001;
font_rom[469] <= 8'b00100000;
font_rom[470] <= 8'b00000001;
font_rom[471] <= 8'b01100000;
font_rom[472] <= 8'b00000011;
font_rom[473] <= 8'b01100000;
font_rom[474] <= 8'b00000011;
font_rom[475] <= 8'b00000000;
font_rom[476] <= 8'b00000000;
font_rom[477] <= 8'b00000000;
font_rom[478] <= 8'b00000000;
font_rom[479] <= 8'b00000000;
//ASCII 0x0F ' '
font_rom[480] <= 8'b00000000;
font_rom[481] <= 8'b00000000;
font_rom[482] <= 8'b00000000;
font_rom[483] <= 8'b00000000;
font_rom[484] <= 8'b00000000;
font_rom[485] <= 8'b00000000;
font_rom[486] <= 8'b00000000;
font_rom[487] <= 8'b00000000;
font_rom[488] <= 8'b00000000;
font_rom[489] <= 8'b00000000;
font_rom[490] <= 8'b00000010;
font_rom[491] <= 8'b10100000;
font_rom[492] <= 8'b00000010;
font_rom[493] <= 8'b10100000;
font_rom[494] <= 8'b00000001;
font_rom[495] <= 8'b01000000;
font_rom[496] <= 8'b00000001;
font_rom[497] <= 8'b01000000;
font_rom[498] <= 8'b00000011;
font_rom[499] <= 8'b01100000;
font_rom[500] <= 8'b00000001;
font_rom[501] <= 8'b01000000;
font_rom[502] <= 8'b00000001;
font_rom[503] <= 8'b01000000;
font_rom[504] <= 8'b00000010;
font_rom[505] <= 8'b10100000;
font_rom[506] <= 8'b00000010;
font_rom[507] <= 8'b10100000;
font_rom[508] <= 8'b00000000;
font_rom[509] <= 8'b00000000;
font_rom[510] <= 8'b00000000;
font_rom[511] <= 8'b00000000;
//ASCII 0x10 ' '
font_rom[512] <= 8'b00000000;
font_rom[513] <= 8'b00000000;
font_rom[514] <= 8'b00000000;
font_rom[515] <= 8'b00000000;
font_rom[516] <= 8'b00000000;
font_rom[517] <= 8'b00000000;
font_rom[518] <= 8'b00000000;
font_rom[519] <= 8'b00000000;
font_rom[520] <= 8'b00000000;
font_rom[521] <= 8'b10000000;
font_rom[522] <= 8'b00000000;
font_rom[523] <= 8'b10000000;
font_rom[524] <= 8'b00000000;
font_rom[525] <= 8'b10000000;
font_rom[526] <= 8'b00000000;
font_rom[527] <= 8'b10000000;
font_rom[528] <= 8'b00000000;
font_rom[529] <= 8'b10000000;
font_rom[530] <= 8'b00000000;
font_rom[531] <= 8'b10000000;
font_rom[532] <= 8'b00000111;
font_rom[533] <= 8'b11100000;
font_rom[534] <= 8'b00000000;
font_rom[535] <= 8'b10000000;
font_rom[536] <= 8'b00000000;
font_rom[537] <= 8'b10000000;
font_rom[538] <= 8'b00000000;
font_rom[539] <= 8'b10000000;
font_rom[540] <= 8'b00000000;
font_rom[541] <= 8'b10000000;
font_rom[542] <= 8'b00000000;
font_rom[543] <= 8'b10000000;
//ASCII 0x11 ' '
font_rom[544] <= 8'b00000000;
font_rom[545] <= 8'b00000000;
font_rom[546] <= 8'b00000000;
font_rom[547] <= 8'b00000000;
font_rom[548] <= 8'b00000000;
font_rom[549] <= 8'b00000000;
font_rom[550] <= 8'b00000000;
font_rom[551] <= 8'b00000000;
font_rom[552] <= 8'b00000000;
font_rom[553] <= 8'b00000000;
font_rom[554] <= 8'b00000000;
font_rom[555] <= 8'b00100000;
font_rom[556] <= 8'b00000000;
font_rom[557] <= 8'b01100000;
font_rom[558] <= 8'b00000000;
font_rom[559] <= 8'b11100000;
font_rom[560] <= 8'b00000001;
font_rom[561] <= 8'b11100000;
font_rom[562] <= 8'b00000011;
font_rom[563] <= 8'b11100000;
font_rom[564] <= 8'b00000001;
font_rom[565] <= 8'b11100000;
font_rom[566] <= 8'b00000000;
font_rom[567] <= 8'b11100000;
font_rom[568] <= 8'b00000000;
font_rom[569] <= 8'b01100000;
font_rom[570] <= 8'b00000000;
font_rom[571] <= 8'b00100000;
font_rom[572] <= 8'b00000000;
font_rom[573] <= 8'b00000000;
font_rom[574] <= 8'b00000000;
font_rom[575] <= 8'b00000000;
//ASCII 0x12 ' '
font_rom[576] <= 8'b00000000;
font_rom[577] <= 8'b00000000;
font_rom[578] <= 8'b00000000;
font_rom[579] <= 8'b00000000;
font_rom[580] <= 8'b00000000;
font_rom[581] <= 8'b00000000;
font_rom[582] <= 8'b00000000;
font_rom[583] <= 8'b00000000;
font_rom[584] <= 8'b00000000;
font_rom[585] <= 8'b10000000;
font_rom[586] <= 8'b00000001;
font_rom[587] <= 8'b11000000;
font_rom[588] <= 8'b00000000;
font_rom[589] <= 8'b10000000;
font_rom[590] <= 8'b00000000;
font_rom[591] <= 8'b10000000;
font_rom[592] <= 8'b00000000;
font_rom[593] <= 8'b10000000;
font_rom[594] <= 8'b00000000;
font_rom[595] <= 8'b10000000;
font_rom[596] <= 8'b00000000;
font_rom[597] <= 8'b10000000;
font_rom[598] <= 8'b00000000;
font_rom[599] <= 8'b10000000;
font_rom[600] <= 8'b00000001;
font_rom[601] <= 8'b11000000;
font_rom[602] <= 8'b00000000;
font_rom[603] <= 8'b10000000;
font_rom[604] <= 8'b00000000;
font_rom[605] <= 8'b00000000;
font_rom[606] <= 8'b00000000;
font_rom[607] <= 8'b00000000;
//ASCII 0x13 ' '
font_rom[608] <= 8'b00000000;
font_rom[609] <= 8'b00000000;
font_rom[610] <= 8'b00000000;
font_rom[611] <= 8'b00000000;
font_rom[612] <= 8'b00000000;
font_rom[613] <= 8'b00000000;
font_rom[614] <= 8'b00000000;
font_rom[615] <= 8'b00000000;
font_rom[616] <= 8'b00000001;
font_rom[617] <= 8'b01000000;
font_rom[618] <= 8'b00000001;
font_rom[619] <= 8'b01000000;
font_rom[620] <= 8'b00000001;
font_rom[621] <= 8'b01000000;
font_rom[622] <= 8'b00000001;
font_rom[623] <= 8'b01000000;
font_rom[624] <= 8'b00000001;
font_rom[625] <= 8'b01000000;
font_rom[626] <= 8'b00000001;
font_rom[627] <= 8'b01000000;
font_rom[628] <= 8'b00000001;
font_rom[629] <= 8'b01000000;
font_rom[630] <= 8'b00000000;
font_rom[631] <= 8'b00000000;
font_rom[632] <= 8'b00000001;
font_rom[633] <= 8'b01000000;
font_rom[634] <= 8'b00000001;
font_rom[635] <= 8'b01000000;
font_rom[636] <= 8'b00000000;
font_rom[637] <= 8'b00000000;
font_rom[638] <= 8'b00000000;
font_rom[639] <= 8'b00000000;
//ASCII 0x14 ' '
font_rom[640] <= 8'b00000000;
font_rom[641] <= 8'b00000000;
font_rom[642] <= 8'b00000000;
font_rom[643] <= 8'b00000000;
font_rom[644] <= 8'b00000000;
font_rom[645] <= 8'b00000000;
font_rom[646] <= 8'b00000000;
font_rom[647] <= 8'b00000000;
font_rom[648] <= 8'b00000001;
font_rom[649] <= 8'b11100000;
font_rom[650] <= 8'b00000010;
font_rom[651] <= 8'b10100000;
font_rom[652] <= 8'b00000010;
font_rom[653] <= 8'b10100000;
font_rom[654] <= 8'b00000010;
font_rom[655] <= 8'b10100000;
font_rom[656] <= 8'b00000001;
font_rom[657] <= 8'b10100000;
font_rom[658] <= 8'b00000000;
font_rom[659] <= 8'b10100000;
font_rom[660] <= 8'b00000000;
font_rom[661] <= 8'b10100000;
font_rom[662] <= 8'b00000000;
font_rom[663] <= 8'b10100000;
font_rom[664] <= 8'b00000000;
font_rom[665] <= 8'b10100000;
font_rom[666] <= 8'b00000000;
font_rom[667] <= 8'b10100000;
font_rom[668] <= 8'b00000000;
font_rom[669] <= 8'b00000000;
font_rom[670] <= 8'b00000000;
font_rom[671] <= 8'b00000000;
//ASCII 0x15 ' '
font_rom[672] <= 8'b00000000;
font_rom[673] <= 8'b00000000;
font_rom[674] <= 8'b00000000;
font_rom[675] <= 8'b00000000;
font_rom[676] <= 8'b00000000;
font_rom[677] <= 8'b00000000;
font_rom[678] <= 8'b00000000;
font_rom[679] <= 8'b00000000;
font_rom[680] <= 8'b00000000;
font_rom[681] <= 8'b10000000;
font_rom[682] <= 8'b00000000;
font_rom[683] <= 8'b10000000;
font_rom[684] <= 8'b00000000;
font_rom[685] <= 8'b10000000;
font_rom[686] <= 8'b00000000;
font_rom[687] <= 8'b10000000;
font_rom[688] <= 8'b00000000;
font_rom[689] <= 8'b10000000;
font_rom[690] <= 8'b00000000;
font_rom[691] <= 8'b10000000;
font_rom[692] <= 8'b00000111;
font_rom[693] <= 8'b11100000;
font_rom[694] <= 8'b00000000;
font_rom[695] <= 8'b00000000;
font_rom[696] <= 8'b00000000;
font_rom[697] <= 8'b00000000;
font_rom[698] <= 8'b00000000;
font_rom[699] <= 8'b00000000;
font_rom[700] <= 8'b00000000;
font_rom[701] <= 8'b00000000;
font_rom[702] <= 8'b00000000;
font_rom[703] <= 8'b00000000;
//ASCII 0x16 ' '
font_rom[704] <= 8'b00000000;
font_rom[705] <= 8'b00000000;
font_rom[706] <= 8'b00000000;
font_rom[707] <= 8'b00000000;
font_rom[708] <= 8'b00000000;
font_rom[709] <= 8'b00000000;
font_rom[710] <= 8'b00000000;
font_rom[711] <= 8'b00000000;
font_rom[712] <= 8'b00000000;
font_rom[713] <= 8'b00000000;
font_rom[714] <= 8'b00000000;
font_rom[715] <= 8'b00000000;
font_rom[716] <= 8'b00000000;
font_rom[717] <= 8'b00000000;
font_rom[718] <= 8'b00000000;
font_rom[719] <= 8'b00000000;
font_rom[720] <= 8'b00000000;
font_rom[721] <= 8'b00000000;
font_rom[722] <= 8'b00000000;
font_rom[723] <= 8'b00000000;
font_rom[724] <= 8'b00000111;
font_rom[725] <= 8'b11100000;
font_rom[726] <= 8'b00000000;
font_rom[727] <= 8'b10000000;
font_rom[728] <= 8'b00000000;
font_rom[729] <= 8'b10000000;
font_rom[730] <= 8'b00000000;
font_rom[731] <= 8'b10000000;
font_rom[732] <= 8'b00000000;
font_rom[733] <= 8'b10000000;
font_rom[734] <= 8'b00000000;
font_rom[735] <= 8'b10000000;
//ASCII 0x17 ' '
font_rom[736] <= 8'b00000000;
font_rom[737] <= 8'b00000000;
font_rom[738] <= 8'b00000000;
font_rom[739] <= 8'b00000000;
font_rom[740] <= 8'b00000000;
font_rom[741] <= 8'b00000000;
font_rom[742] <= 8'b00000000;
font_rom[743] <= 8'b00000000;
font_rom[744] <= 8'b00000000;
font_rom[745] <= 8'b10000000;
font_rom[746] <= 8'b00000000;
font_rom[747] <= 8'b10000000;
font_rom[748] <= 8'b00000000;
font_rom[749] <= 8'b10000000;
font_rom[750] <= 8'b00000000;
font_rom[751] <= 8'b10000000;
font_rom[752] <= 8'b00000000;
font_rom[753] <= 8'b10000000;
font_rom[754] <= 8'b00000000;
font_rom[755] <= 8'b10000000;
font_rom[756] <= 8'b00000111;
font_rom[757] <= 8'b10000000;
font_rom[758] <= 8'b00000000;
font_rom[759] <= 8'b10000000;
font_rom[760] <= 8'b00000000;
font_rom[761] <= 8'b10000000;
font_rom[762] <= 8'b00000000;
font_rom[763] <= 8'b10000000;
font_rom[764] <= 8'b00000000;
font_rom[765] <= 8'b10000000;
font_rom[766] <= 8'b00000000;
font_rom[767] <= 8'b10000000;
//ASCII 0x18 ' '
font_rom[768] <= 8'b00000000;
font_rom[769] <= 8'b00000000;
font_rom[770] <= 8'b00000000;
font_rom[771] <= 8'b00000000;
font_rom[772] <= 8'b00000000;
font_rom[773] <= 8'b00000000;
font_rom[774] <= 8'b00000000;
font_rom[775] <= 8'b00000000;
font_rom[776] <= 8'b00000000;
font_rom[777] <= 8'b10000000;
font_rom[778] <= 8'b00000001;
font_rom[779] <= 8'b11000000;
font_rom[780] <= 8'b00000000;
font_rom[781] <= 8'b10000000;
font_rom[782] <= 8'b00000000;
font_rom[783] <= 8'b10000000;
font_rom[784] <= 8'b00000000;
font_rom[785] <= 8'b10000000;
font_rom[786] <= 8'b00000000;
font_rom[787] <= 8'b10000000;
font_rom[788] <= 8'b00000000;
font_rom[789] <= 8'b10000000;
font_rom[790] <= 8'b00000000;
font_rom[791] <= 8'b10000000;
font_rom[792] <= 8'b00000000;
font_rom[793] <= 8'b10000000;
font_rom[794] <= 8'b00000000;
font_rom[795] <= 8'b10000000;
font_rom[796] <= 8'b00000000;
font_rom[797] <= 8'b00000000;
font_rom[798] <= 8'b00000000;
font_rom[799] <= 8'b00000000;
//ASCII 0x19 ' '
font_rom[800] <= 8'b00000000;
font_rom[801] <= 8'b00000000;
font_rom[802] <= 8'b00000000;
font_rom[803] <= 8'b00000000;
font_rom[804] <= 8'b00000000;
font_rom[805] <= 8'b00000000;
font_rom[806] <= 8'b00000000;
font_rom[807] <= 8'b00000000;
font_rom[808] <= 8'b00000000;
font_rom[809] <= 8'b10000000;
font_rom[810] <= 8'b00000000;
font_rom[811] <= 8'b10000000;
font_rom[812] <= 8'b00000000;
font_rom[813] <= 8'b10000000;
font_rom[814] <= 8'b00000000;
font_rom[815] <= 8'b10000000;
font_rom[816] <= 8'b00000000;
font_rom[817] <= 8'b10000000;
font_rom[818] <= 8'b00000000;
font_rom[819] <= 8'b10000000;
font_rom[820] <= 8'b00000000;
font_rom[821] <= 8'b11100000;
font_rom[822] <= 8'b00000000;
font_rom[823] <= 8'b10000000;
font_rom[824] <= 8'b00000000;
font_rom[825] <= 8'b10000000;
font_rom[826] <= 8'b00000000;
font_rom[827] <= 8'b10000000;
font_rom[828] <= 8'b00000000;
font_rom[829] <= 8'b10000000;
font_rom[830] <= 8'b00000000;
font_rom[831] <= 8'b10000000;
//ASCII 0x1A ' '
font_rom[832] <= 8'b00000000;
font_rom[833] <= 8'b00000000;
font_rom[834] <= 8'b00000000;
font_rom[835] <= 8'b00000000;
font_rom[836] <= 8'b00000000;
font_rom[837] <= 8'b00000000;
font_rom[838] <= 8'b00000000;
font_rom[839] <= 8'b00000000;
font_rom[840] <= 8'b00000000;
font_rom[841] <= 8'b00000000;
font_rom[842] <= 8'b00000000;
font_rom[843] <= 8'b00000000;
font_rom[844] <= 8'b00000000;
font_rom[845] <= 8'b00000000;
font_rom[846] <= 8'b00000000;
font_rom[847] <= 8'b00000000;
font_rom[848] <= 8'b00000000;
font_rom[849] <= 8'b01000000;
font_rom[850] <= 8'b00000011;
font_rom[851] <= 8'b11100000;
font_rom[852] <= 8'b00000000;
font_rom[853] <= 8'b01000000;
font_rom[854] <= 8'b00000000;
font_rom[855] <= 8'b00000000;
font_rom[856] <= 8'b00000000;
font_rom[857] <= 8'b00000000;
font_rom[858] <= 8'b00000000;
font_rom[859] <= 8'b00000000;
font_rom[860] <= 8'b00000000;
font_rom[861] <= 8'b00000000;
font_rom[862] <= 8'b00000000;
font_rom[863] <= 8'b00000000;
//ASCII 0x1B ' '
font_rom[864] <= 8'b00000000;
font_rom[865] <= 8'b00000000;
font_rom[866] <= 8'b00000000;
font_rom[867] <= 8'b00000000;
font_rom[868] <= 8'b00000000;
font_rom[869] <= 8'b00000000;
font_rom[870] <= 8'b00000000;
font_rom[871] <= 8'b00000000;
font_rom[872] <= 8'b00000000;
font_rom[873] <= 8'b00000000;
font_rom[874] <= 8'b00000000;
font_rom[875] <= 8'b00000000;
font_rom[876] <= 8'b00000000;
font_rom[877] <= 8'b00000000;
font_rom[878] <= 8'b00000000;
font_rom[879] <= 8'b00000000;
font_rom[880] <= 8'b00000001;
font_rom[881] <= 8'b00000000;
font_rom[882] <= 8'b00000011;
font_rom[883] <= 8'b11100000;
font_rom[884] <= 8'b00000001;
font_rom[885] <= 8'b00000000;
font_rom[886] <= 8'b00000000;
font_rom[887] <= 8'b00000000;
font_rom[888] <= 8'b00000000;
font_rom[889] <= 8'b00000000;
font_rom[890] <= 8'b00000000;
font_rom[891] <= 8'b00000000;
font_rom[892] <= 8'b00000000;
font_rom[893] <= 8'b00000000;
font_rom[894] <= 8'b00000000;
font_rom[895] <= 8'b00000000;
//ASCII 0x1C ' '
font_rom[896] <= 8'b00000000;
font_rom[897] <= 8'b00000000;
font_rom[898] <= 8'b00000000;
font_rom[899] <= 8'b00000000;
font_rom[900] <= 8'b00000000;
font_rom[901] <= 8'b00000000;
font_rom[902] <= 8'b00000000;
font_rom[903] <= 8'b00000000;
font_rom[904] <= 8'b00000000;
font_rom[905] <= 8'b00000000;
font_rom[906] <= 8'b00000000;
font_rom[907] <= 8'b00000000;
font_rom[908] <= 8'b00000000;
font_rom[909] <= 8'b00000000;
font_rom[910] <= 8'b00000000;
font_rom[911] <= 8'b00000000;
font_rom[912] <= 8'b00000000;
font_rom[913] <= 8'b00000000;
font_rom[914] <= 8'b00000000;
font_rom[915] <= 8'b00000000;
font_rom[916] <= 8'b00000000;
font_rom[917] <= 8'b00000000;
font_rom[918] <= 8'b00000000;
font_rom[919] <= 8'b00000000;
font_rom[920] <= 8'b00000000;
font_rom[921] <= 8'b00000000;
font_rom[922] <= 8'b00000000;
font_rom[923] <= 8'b00000000;
font_rom[924] <= 8'b00000000;
font_rom[925] <= 8'b00000000;
font_rom[926] <= 8'b00000000;
font_rom[927] <= 8'b00000000;
//ASCII 0x1D ' '
font_rom[928] <= 8'b00000000;
font_rom[929] <= 8'b00000000;
font_rom[930] <= 8'b00000000;
font_rom[931] <= 8'b00000000;
font_rom[932] <= 8'b00000000;
font_rom[933] <= 8'b00000000;
font_rom[934] <= 8'b00000000;
font_rom[935] <= 8'b00000000;
font_rom[936] <= 8'b00000000;
font_rom[937] <= 8'b00000000;
font_rom[938] <= 8'b00000000;
font_rom[939] <= 8'b00000000;
font_rom[940] <= 8'b00000000;
font_rom[941] <= 8'b00000000;
font_rom[942] <= 8'b00000000;
font_rom[943] <= 8'b00000000;
font_rom[944] <= 8'b00000000;
font_rom[945] <= 8'b00000000;
font_rom[946] <= 8'b00000000;
font_rom[947] <= 8'b00000000;
font_rom[948] <= 8'b00000000;
font_rom[949] <= 8'b00000000;
font_rom[950] <= 8'b00000000;
font_rom[951] <= 8'b00000000;
font_rom[952] <= 8'b00000000;
font_rom[953] <= 8'b00000000;
font_rom[954] <= 8'b00000000;
font_rom[955] <= 8'b00000000;
font_rom[956] <= 8'b00000000;
font_rom[957] <= 8'b00000000;
font_rom[958] <= 8'b00000000;
font_rom[959] <= 8'b00000000;
//ASCII 0x1E ' '
font_rom[960] <= 8'b00000000;
font_rom[961] <= 8'b00000000;
font_rom[962] <= 8'b00000000;
font_rom[963] <= 8'b00000000;
font_rom[964] <= 8'b00000000;
font_rom[965] <= 8'b00000000;
font_rom[966] <= 8'b00000000;
font_rom[967] <= 8'b00000000;
font_rom[968] <= 8'b00000000;
font_rom[969] <= 8'b00000000;
font_rom[970] <= 8'b00000000;
font_rom[971] <= 8'b00000000;
font_rom[972] <= 8'b00000000;
font_rom[973] <= 8'b00000000;
font_rom[974] <= 8'b00000000;
font_rom[975] <= 8'b00000000;
font_rom[976] <= 8'b00000000;
font_rom[977] <= 8'b00000000;
font_rom[978] <= 8'b00000000;
font_rom[979] <= 8'b00000000;
font_rom[980] <= 8'b00000000;
font_rom[981] <= 8'b00000000;
font_rom[982] <= 8'b00000000;
font_rom[983] <= 8'b00000000;
font_rom[984] <= 8'b00000000;
font_rom[985] <= 8'b00000000;
font_rom[986] <= 8'b00000000;
font_rom[987] <= 8'b00000000;
font_rom[988] <= 8'b00000000;
font_rom[989] <= 8'b00000000;
font_rom[990] <= 8'b00000000;
font_rom[991] <= 8'b00000000;
//ASCII 0x1F ' '
font_rom[992] <= 8'b00000000;
font_rom[993] <= 8'b00000000;
font_rom[994] <= 8'b00000000;
font_rom[995] <= 8'b00000000;
font_rom[996] <= 8'b00000000;
font_rom[997] <= 8'b00000000;
font_rom[998] <= 8'b00000000;
font_rom[999] <= 8'b00000000;
font_rom[1000] <= 8'b00000000;
font_rom[1001] <= 8'b00000000;
font_rom[1002] <= 8'b00000000;
font_rom[1003] <= 8'b00000000;
font_rom[1004] <= 8'b00000000;
font_rom[1005] <= 8'b00000000;
font_rom[1006] <= 8'b00000000;
font_rom[1007] <= 8'b00000000;
font_rom[1008] <= 8'b00000000;
font_rom[1009] <= 8'b00000000;
font_rom[1010] <= 8'b00000000;
font_rom[1011] <= 8'b00000000;
font_rom[1012] <= 8'b00000000;
font_rom[1013] <= 8'b00000000;
font_rom[1014] <= 8'b00000000;
font_rom[1015] <= 8'b00000000;
font_rom[1016] <= 8'b00000000;
font_rom[1017] <= 8'b00000000;
font_rom[1018] <= 8'b00000000;
font_rom[1019] <= 8'b00000000;
font_rom[1020] <= 8'b00000000;
font_rom[1021] <= 8'b00000000;
font_rom[1022] <= 8'b00000000;
font_rom[1023] <= 8'b00000000;
//ASCII 0x20 ' '
font_rom[1024] <= 8'b00000000;
font_rom[1025] <= 8'b00000000;
font_rom[1026] <= 8'b00000000;
font_rom[1027] <= 8'b00000000;
font_rom[1028] <= 8'b00000000;
font_rom[1029] <= 8'b00000000;
font_rom[1030] <= 8'b00000000;
font_rom[1031] <= 8'b00000000;
font_rom[1032] <= 8'b00000000;
font_rom[1033] <= 8'b00000000;
font_rom[1034] <= 8'b00000000;
font_rom[1035] <= 8'b00000000;
font_rom[1036] <= 8'b00000000;
font_rom[1037] <= 8'b00000000;
font_rom[1038] <= 8'b00000000;
font_rom[1039] <= 8'b00000000;
font_rom[1040] <= 8'b00000000;
font_rom[1041] <= 8'b00000000;
font_rom[1042] <= 8'b00000000;
font_rom[1043] <= 8'b00000000;
font_rom[1044] <= 8'b00000000;
font_rom[1045] <= 8'b00000000;
font_rom[1046] <= 8'b00000000;
font_rom[1047] <= 8'b00000000;
font_rom[1048] <= 8'b00000000;
font_rom[1049] <= 8'b00000000;
font_rom[1050] <= 8'b00000000;
font_rom[1051] <= 8'b00000000;
font_rom[1052] <= 8'b00000000;
font_rom[1053] <= 8'b00000000;
font_rom[1054] <= 8'b00000000;
font_rom[1055] <= 8'b00000000;
//ASCII 0x21 '!'
font_rom[1056] <= 8'b00000000;
font_rom[1057] <= 8'b00000000;
font_rom[1058] <= 8'b00000000;
font_rom[1059] <= 8'b00000000;
font_rom[1060] <= 8'b00000000;
font_rom[1061] <= 8'b00000000;
font_rom[1062] <= 8'b00000000;
font_rom[1063] <= 8'b00000000;
font_rom[1064] <= 8'b00000011;
font_rom[1065] <= 8'b00000000;
font_rom[1066] <= 8'b00000011;
font_rom[1067] <= 8'b00000000;
font_rom[1068] <= 8'b00000011;
font_rom[1069] <= 8'b00000000;
font_rom[1070] <= 8'b00000011;
font_rom[1071] <= 8'b00000000;
font_rom[1072] <= 8'b00000011;
font_rom[1073] <= 8'b00000000;
font_rom[1074] <= 8'b00000011;
font_rom[1075] <= 8'b00000000;
font_rom[1076] <= 8'b00000011;
font_rom[1077] <= 8'b00000000;
font_rom[1078] <= 8'b00000000;
font_rom[1079] <= 8'b00000000;
font_rom[1080] <= 8'b00000011;
font_rom[1081] <= 8'b00000000;
font_rom[1082] <= 8'b00000000;
font_rom[1083] <= 8'b00000000;
font_rom[1084] <= 8'b00000000;
font_rom[1085] <= 8'b00000000;
font_rom[1086] <= 8'b00000000;
font_rom[1087] <= 8'b00000000;
//ASCII 0x22 '"'
font_rom[1088] <= 8'b00000000;
font_rom[1089] <= 8'b00000000;
font_rom[1090] <= 8'b00000000;
font_rom[1091] <= 8'b00000000;
font_rom[1092] <= 8'b00000000;
font_rom[1093] <= 8'b00000000;
font_rom[1094] <= 8'b00000000;
font_rom[1095] <= 8'b00000000;
font_rom[1096] <= 8'b00000000;
font_rom[1097] <= 8'b00000000;
font_rom[1098] <= 8'b00000011;
font_rom[1099] <= 8'b11000000;
font_rom[1100] <= 8'b00000011;
font_rom[1101] <= 8'b11000000;
font_rom[1102] <= 8'b00000011;
font_rom[1103] <= 8'b11000000;
font_rom[1104] <= 8'b00000000;
font_rom[1105] <= 8'b00000000;
font_rom[1106] <= 8'b00000000;
font_rom[1107] <= 8'b00000000;
font_rom[1108] <= 8'b00000000;
font_rom[1109] <= 8'b00000000;
font_rom[1110] <= 8'b00000000;
font_rom[1111] <= 8'b00000000;
font_rom[1112] <= 8'b00000000;
font_rom[1113] <= 8'b00000000;
font_rom[1114] <= 8'b00000000;
font_rom[1115] <= 8'b00000000;
font_rom[1116] <= 8'b00000000;
font_rom[1117] <= 8'b00000000;
font_rom[1118] <= 8'b00000000;
font_rom[1119] <= 8'b00000000;
//ASCII 0x23 '#'
font_rom[1120] <= 8'b00000000;
font_rom[1121] <= 8'b00000000;
font_rom[1122] <= 8'b00000000;
font_rom[1123] <= 8'b00000000;
font_rom[1124] <= 8'b00000000;
font_rom[1125] <= 8'b00000000;
font_rom[1126] <= 8'b00000000;
font_rom[1127] <= 8'b00000000;
font_rom[1128] <= 8'b00000000;
font_rom[1129] <= 8'b00000000;
font_rom[1130] <= 8'b00000001;
font_rom[1131] <= 8'b00110000;
font_rom[1132] <= 8'b00000011;
font_rom[1133] <= 8'b00110000;
font_rom[1134] <= 8'b00001111;
font_rom[1135] <= 8'b11111000;
font_rom[1136] <= 8'b00000011;
font_rom[1137] <= 8'b01100000;
font_rom[1138] <= 8'b00000110;
font_rom[1139] <= 8'b01100000;
font_rom[1140] <= 8'b00011111;
font_rom[1141] <= 8'b11111000;
font_rom[1142] <= 8'b00000110;
font_rom[1143] <= 8'b11000000;
font_rom[1144] <= 8'b00001100;
font_rom[1145] <= 8'b11000000;
font_rom[1146] <= 8'b00000000;
font_rom[1147] <= 8'b00000000;
font_rom[1148] <= 8'b00000000;
font_rom[1149] <= 8'b00000000;
font_rom[1150] <= 8'b00000000;
font_rom[1151] <= 8'b00000000;
//ASCII 0x24 '$'
font_rom[1152] <= 8'b00000000;
font_rom[1153] <= 8'b00000000;
font_rom[1154] <= 8'b00000000;
font_rom[1155] <= 8'b00000000;
font_rom[1156] <= 8'b00000000;
font_rom[1157] <= 8'b00000000;
font_rom[1158] <= 8'b00000000;
font_rom[1159] <= 8'b00000000;
font_rom[1160] <= 8'b00000011;
font_rom[1161] <= 8'b00000000;
font_rom[1162] <= 8'b00000111;
font_rom[1163] <= 8'b11100000;
font_rom[1164] <= 8'b00001111;
font_rom[1165] <= 8'b00000000;
font_rom[1166] <= 8'b00001111;
font_rom[1167] <= 8'b00000000;
font_rom[1168] <= 8'b00000111;
font_rom[1169] <= 8'b11000000;
font_rom[1170] <= 8'b00000011;
font_rom[1171] <= 8'b01100000;
font_rom[1172] <= 8'b00000011;
font_rom[1173] <= 8'b01100000;
font_rom[1174] <= 8'b00000011;
font_rom[1175] <= 8'b11100000;
font_rom[1176] <= 8'b00001111;
font_rom[1177] <= 8'b11000000;
font_rom[1178] <= 8'b00000011;
font_rom[1179] <= 8'b00000000;
font_rom[1180] <= 8'b00000011;
font_rom[1181] <= 8'b00000000;
font_rom[1182] <= 8'b00000000;
font_rom[1183] <= 8'b00000000;
//ASCII 0x25 '%'
font_rom[1184] <= 8'b00000000;
font_rom[1185] <= 8'b00000000;
font_rom[1186] <= 8'b00000000;
font_rom[1187] <= 8'b00000000;
font_rom[1188] <= 8'b00000000;
font_rom[1189] <= 8'b00000000;
font_rom[1190] <= 8'b00000000;
font_rom[1191] <= 8'b00000000;
font_rom[1192] <= 8'b00000000;
font_rom[1193] <= 8'b01100000;
font_rom[1194] <= 8'b00000111;
font_rom[1195] <= 8'b01000000;
font_rom[1196] <= 8'b00001111;
font_rom[1197] <= 8'b11000000;
font_rom[1198] <= 8'b00001111;
font_rom[1199] <= 8'b11000000;
font_rom[1200] <= 8'b00000111;
font_rom[1201] <= 8'b10000000;
font_rom[1202] <= 8'b00000001;
font_rom[1203] <= 8'b11110000;
font_rom[1204] <= 8'b00000011;
font_rom[1205] <= 8'b11011000;
font_rom[1206] <= 8'b00000011;
font_rom[1207] <= 8'b11011000;
font_rom[1208] <= 8'b00000110;
font_rom[1209] <= 8'b01110000;
font_rom[1210] <= 8'b00000000;
font_rom[1211] <= 8'b00000000;
font_rom[1212] <= 8'b00000000;
font_rom[1213] <= 8'b00000000;
font_rom[1214] <= 8'b00000000;
font_rom[1215] <= 8'b00000000;
//ASCII 0x26 '&'
font_rom[1216] <= 8'b00000000;
font_rom[1217] <= 8'b00000000;
font_rom[1218] <= 8'b00000000;
font_rom[1219] <= 8'b00000000;
font_rom[1220] <= 8'b00000000;
font_rom[1221] <= 8'b00000000;
font_rom[1222] <= 8'b00000000;
font_rom[1223] <= 8'b00000000;
font_rom[1224] <= 8'b00000000;
font_rom[1225] <= 8'b00000000;
font_rom[1226] <= 8'b00000011;
font_rom[1227] <= 8'b10000000;
font_rom[1228] <= 8'b00000011;
font_rom[1229] <= 8'b10000000;
font_rom[1230] <= 8'b00000011;
font_rom[1231] <= 8'b10000000;
font_rom[1232] <= 8'b00000111;
font_rom[1233] <= 8'b01100000;
font_rom[1234] <= 8'b00001101;
font_rom[1235] <= 8'b11100000;
font_rom[1236] <= 8'b00001100;
font_rom[1237] <= 8'b11000000;
font_rom[1238] <= 8'b00001100;
font_rom[1239] <= 8'b11000000;
font_rom[1240] <= 8'b00000111;
font_rom[1241] <= 8'b11100000;
font_rom[1242] <= 8'b00000000;
font_rom[1243] <= 8'b00000000;
font_rom[1244] <= 8'b00000000;
font_rom[1245] <= 8'b00000000;
font_rom[1246] <= 8'b00000000;
font_rom[1247] <= 8'b00000000;
//ASCII 0x27 '''
font_rom[1248] <= 8'b00000000;
font_rom[1249] <= 8'b00000000;
font_rom[1250] <= 8'b00000000;
font_rom[1251] <= 8'b00000000;
font_rom[1252] <= 8'b00000000;
font_rom[1253] <= 8'b00000000;
font_rom[1254] <= 8'b00000000;
font_rom[1255] <= 8'b00000000;
font_rom[1256] <= 8'b00000000;
font_rom[1257] <= 8'b00000000;
font_rom[1258] <= 8'b00000001;
font_rom[1259] <= 8'b10000000;
font_rom[1260] <= 8'b00000001;
font_rom[1261] <= 8'b10000000;
font_rom[1262] <= 8'b00000001;
font_rom[1263] <= 8'b10000000;
font_rom[1264] <= 8'b00000000;
font_rom[1265] <= 8'b00000000;
font_rom[1266] <= 8'b00000000;
font_rom[1267] <= 8'b00000000;
font_rom[1268] <= 8'b00000000;
font_rom[1269] <= 8'b00000000;
font_rom[1270] <= 8'b00000000;
font_rom[1271] <= 8'b00000000;
font_rom[1272] <= 8'b00000000;
font_rom[1273] <= 8'b00000000;
font_rom[1274] <= 8'b00000000;
font_rom[1275] <= 8'b00000000;
font_rom[1276] <= 8'b00000000;
font_rom[1277] <= 8'b00000000;
font_rom[1278] <= 8'b00000000;
font_rom[1279] <= 8'b00000000;
//ASCII 0x28 '('
font_rom[1280] <= 8'b00000000;
font_rom[1281] <= 8'b00000000;
font_rom[1282] <= 8'b00000000;
font_rom[1283] <= 8'b00000000;
font_rom[1284] <= 8'b00000000;
font_rom[1285] <= 8'b00000000;
font_rom[1286] <= 8'b00000000;
font_rom[1287] <= 8'b00000000;
font_rom[1288] <= 8'b00000000;
font_rom[1289] <= 8'b11000000;
font_rom[1290] <= 8'b00000001;
font_rom[1291] <= 8'b10000000;
font_rom[1292] <= 8'b00000011;
font_rom[1293] <= 8'b00000000;
font_rom[1294] <= 8'b00000011;
font_rom[1295] <= 8'b00000000;
font_rom[1296] <= 8'b00000011;
font_rom[1297] <= 8'b00000000;
font_rom[1298] <= 8'b00000011;
font_rom[1299] <= 8'b00000000;
font_rom[1300] <= 8'b00000011;
font_rom[1301] <= 8'b00000000;
font_rom[1302] <= 8'b00000011;
font_rom[1303] <= 8'b00000000;
font_rom[1304] <= 8'b00000011;
font_rom[1305] <= 8'b00000000;
font_rom[1306] <= 8'b00000001;
font_rom[1307] <= 8'b10000000;
font_rom[1308] <= 8'b00000000;
font_rom[1309] <= 8'b11000000;
font_rom[1310] <= 8'b00000000;
font_rom[1311] <= 8'b00000000;
//ASCII 0x29 ')'
font_rom[1312] <= 8'b00000000;
font_rom[1313] <= 8'b00000000;
font_rom[1314] <= 8'b00000000;
font_rom[1315] <= 8'b00000000;
font_rom[1316] <= 8'b00000000;
font_rom[1317] <= 8'b00000000;
font_rom[1318] <= 8'b00000000;
font_rom[1319] <= 8'b00000000;
font_rom[1320] <= 8'b00000011;
font_rom[1321] <= 8'b00000000;
font_rom[1322] <= 8'b00000011;
font_rom[1323] <= 8'b10000000;
font_rom[1324] <= 8'b00000001;
font_rom[1325] <= 8'b10000000;
font_rom[1326] <= 8'b00000001;
font_rom[1327] <= 8'b10000000;
font_rom[1328] <= 8'b00000000;
font_rom[1329] <= 8'b11000000;
font_rom[1330] <= 8'b00000000;
font_rom[1331] <= 8'b11000000;
font_rom[1332] <= 8'b00000000;
font_rom[1333] <= 8'b11000000;
font_rom[1334] <= 8'b00000000;
font_rom[1335] <= 8'b10000000;
font_rom[1336] <= 8'b00000001;
font_rom[1337] <= 8'b10000000;
font_rom[1338] <= 8'b00000001;
font_rom[1339] <= 8'b10000000;
font_rom[1340] <= 8'b00000011;
font_rom[1341] <= 8'b00000000;
font_rom[1342] <= 8'b00000000;
font_rom[1343] <= 8'b00000000;
//ASCII 0x2A '*'
font_rom[1344] <= 8'b00000000;
font_rom[1345] <= 8'b00000000;
font_rom[1346] <= 8'b00000000;
font_rom[1347] <= 8'b00000000;
font_rom[1348] <= 8'b00000000;
font_rom[1349] <= 8'b00000000;
font_rom[1350] <= 8'b00000000;
font_rom[1351] <= 8'b00000000;
font_rom[1352] <= 8'b00000000;
font_rom[1353] <= 8'b00000000;
font_rom[1354] <= 8'b00000011;
font_rom[1355] <= 8'b00000000;
font_rom[1356] <= 8'b00000111;
font_rom[1357] <= 8'b11000000;
font_rom[1358] <= 8'b00000011;
font_rom[1359] <= 8'b10000000;
font_rom[1360] <= 8'b00000110;
font_rom[1361] <= 8'b11000000;
font_rom[1362] <= 8'b00000000;
font_rom[1363] <= 8'b00000000;
font_rom[1364] <= 8'b00000000;
font_rom[1365] <= 8'b00000000;
font_rom[1366] <= 8'b00000000;
font_rom[1367] <= 8'b00000000;
font_rom[1368] <= 8'b00000000;
font_rom[1369] <= 8'b00000000;
font_rom[1370] <= 8'b00000000;
font_rom[1371] <= 8'b00000000;
font_rom[1372] <= 8'b00000000;
font_rom[1373] <= 8'b00000000;
font_rom[1374] <= 8'b00000000;
font_rom[1375] <= 8'b00000000;
//ASCII 0x2B '+'
font_rom[1376] <= 8'b00000000;
font_rom[1377] <= 8'b00000000;
font_rom[1378] <= 8'b00000000;
font_rom[1379] <= 8'b00000000;
font_rom[1380] <= 8'b00000000;
font_rom[1381] <= 8'b00000000;
font_rom[1382] <= 8'b00000000;
font_rom[1383] <= 8'b00000000;
font_rom[1384] <= 8'b00000000;
font_rom[1385] <= 8'b00000000;
font_rom[1386] <= 8'b00000000;
font_rom[1387] <= 8'b00000000;
font_rom[1388] <= 8'b00000000;
font_rom[1389] <= 8'b00000000;
font_rom[1390] <= 8'b00000001;
font_rom[1391] <= 8'b10000000;
font_rom[1392] <= 8'b00000001;
font_rom[1393] <= 8'b10000000;
font_rom[1394] <= 8'b00000111;
font_rom[1395] <= 8'b11100000;
font_rom[1396] <= 8'b00000001;
font_rom[1397] <= 8'b10000000;
font_rom[1398] <= 8'b00000001;
font_rom[1399] <= 8'b10000000;
font_rom[1400] <= 8'b00000000;
font_rom[1401] <= 8'b00000000;
font_rom[1402] <= 8'b00000000;
font_rom[1403] <= 8'b00000000;
font_rom[1404] <= 8'b00000000;
font_rom[1405] <= 8'b00000000;
font_rom[1406] <= 8'b00000000;
font_rom[1407] <= 8'b00000000;
//ASCII 0x2C ','
font_rom[1408] <= 8'b00000000;
font_rom[1409] <= 8'b00000000;
font_rom[1410] <= 8'b00000000;
font_rom[1411] <= 8'b00000000;
font_rom[1412] <= 8'b00000000;
font_rom[1413] <= 8'b00000000;
font_rom[1414] <= 8'b00000000;
font_rom[1415] <= 8'b00000000;
font_rom[1416] <= 8'b00000000;
font_rom[1417] <= 8'b00000000;
font_rom[1418] <= 8'b00000000;
font_rom[1419] <= 8'b00000000;
font_rom[1420] <= 8'b00000000;
font_rom[1421] <= 8'b00000000;
font_rom[1422] <= 8'b00000000;
font_rom[1423] <= 8'b00000000;
font_rom[1424] <= 8'b00000000;
font_rom[1425] <= 8'b00000000;
font_rom[1426] <= 8'b00000000;
font_rom[1427] <= 8'b00000000;
font_rom[1428] <= 8'b00000000;
font_rom[1429] <= 8'b00000000;
font_rom[1430] <= 8'b00000000;
font_rom[1431] <= 8'b00000000;
font_rom[1432] <= 8'b00000001;
font_rom[1433] <= 8'b10000000;
font_rom[1434] <= 8'b00000011;
font_rom[1435] <= 8'b00000000;
font_rom[1436] <= 8'b00000000;
font_rom[1437] <= 8'b00000000;
font_rom[1438] <= 8'b00000000;
font_rom[1439] <= 8'b00000000;
//ASCII 0x2D '-'
font_rom[1440] <= 8'b00000000;
font_rom[1441] <= 8'b00000000;
font_rom[1442] <= 8'b00000000;
font_rom[1443] <= 8'b00000000;
font_rom[1444] <= 8'b00000000;
font_rom[1445] <= 8'b00000000;
font_rom[1446] <= 8'b00000000;
font_rom[1447] <= 8'b00000000;
font_rom[1448] <= 8'b00000000;
font_rom[1449] <= 8'b00000000;
font_rom[1450] <= 8'b00000000;
font_rom[1451] <= 8'b00000000;
font_rom[1452] <= 8'b00000000;
font_rom[1453] <= 8'b00000000;
font_rom[1454] <= 8'b00000000;
font_rom[1455] <= 8'b00000000;
font_rom[1456] <= 8'b00000000;
font_rom[1457] <= 8'b00000000;
font_rom[1458] <= 8'b00000000;
font_rom[1459] <= 8'b00000000;
font_rom[1460] <= 8'b00000011;
font_rom[1461] <= 8'b11000000;
font_rom[1462] <= 8'b00000000;
font_rom[1463] <= 8'b00000000;
font_rom[1464] <= 8'b00000000;
font_rom[1465] <= 8'b00000000;
font_rom[1466] <= 8'b00000000;
font_rom[1467] <= 8'b00000000;
font_rom[1468] <= 8'b00000000;
font_rom[1469] <= 8'b00000000;
font_rom[1470] <= 8'b00000000;
font_rom[1471] <= 8'b00000000;
//ASCII 0x2E '.'
font_rom[1472] <= 8'b00000000;
font_rom[1473] <= 8'b00000000;
font_rom[1474] <= 8'b00000000;
font_rom[1475] <= 8'b00000000;
font_rom[1476] <= 8'b00000000;
font_rom[1477] <= 8'b00000000;
font_rom[1478] <= 8'b00000000;
font_rom[1479] <= 8'b00000000;
font_rom[1480] <= 8'b00000000;
font_rom[1481] <= 8'b00000000;
font_rom[1482] <= 8'b00000000;
font_rom[1483] <= 8'b00000000;
font_rom[1484] <= 8'b00000000;
font_rom[1485] <= 8'b00000000;
font_rom[1486] <= 8'b00000000;
font_rom[1487] <= 8'b00000000;
font_rom[1488] <= 8'b00000000;
font_rom[1489] <= 8'b00000000;
font_rom[1490] <= 8'b00000000;
font_rom[1491] <= 8'b00000000;
font_rom[1492] <= 8'b00000000;
font_rom[1493] <= 8'b00000000;
font_rom[1494] <= 8'b00000000;
font_rom[1495] <= 8'b00000000;
font_rom[1496] <= 8'b00000011;
font_rom[1497] <= 8'b00000000;
font_rom[1498] <= 8'b00000000;
font_rom[1499] <= 8'b00000000;
font_rom[1500] <= 8'b00000000;
font_rom[1501] <= 8'b00000000;
font_rom[1502] <= 8'b00000000;
font_rom[1503] <= 8'b00000000;
//ASCII 0x2F '/'
font_rom[1504] <= 8'b00000000;
font_rom[1505] <= 8'b00000000;
font_rom[1506] <= 8'b00000000;
font_rom[1507] <= 8'b00000000;
font_rom[1508] <= 8'b00000000;
font_rom[1509] <= 8'b00000000;
font_rom[1510] <= 8'b00000000;
font_rom[1511] <= 8'b00000000;
font_rom[1512] <= 8'b00000000;
font_rom[1513] <= 8'b11000000;
font_rom[1514] <= 8'b00000000;
font_rom[1515] <= 8'b11000000;
font_rom[1516] <= 8'b00000000;
font_rom[1517] <= 8'b10000000;
font_rom[1518] <= 8'b00000001;
font_rom[1519] <= 8'b10000000;
font_rom[1520] <= 8'b00000001;
font_rom[1521] <= 8'b00000000;
font_rom[1522] <= 8'b00000011;
font_rom[1523] <= 8'b00000000;
font_rom[1524] <= 8'b00000010;
font_rom[1525] <= 8'b00000000;
font_rom[1526] <= 8'b00000110;
font_rom[1527] <= 8'b00000000;
font_rom[1528] <= 8'b00000110;
font_rom[1529] <= 8'b00000000;
font_rom[1530] <= 8'b00000000;
font_rom[1531] <= 8'b00000000;
font_rom[1532] <= 8'b00000000;
font_rom[1533] <= 8'b00000000;
font_rom[1534] <= 8'b00000000;
font_rom[1535] <= 8'b00000000;
//ASCII 0x30 '0'
font_rom[1536] <= 8'b00000000;
font_rom[1537] <= 8'b00000000;
font_rom[1538] <= 8'b00000000;
font_rom[1539] <= 8'b00000000;
font_rom[1540] <= 8'b00000000;
font_rom[1541] <= 8'b00000000;
font_rom[1542] <= 8'b00000000;
font_rom[1543] <= 8'b00000000;
font_rom[1544] <= 8'b00000000;
font_rom[1545] <= 8'b00000000;
font_rom[1546] <= 8'b00000111;
font_rom[1547] <= 8'b11000000;
font_rom[1548] <= 8'b00001100;
font_rom[1549] <= 8'b11000000;
font_rom[1550] <= 8'b00001100;
font_rom[1551] <= 8'b01000000;
font_rom[1552] <= 8'b00001000;
font_rom[1553] <= 8'b01100000;
font_rom[1554] <= 8'b00001000;
font_rom[1555] <= 8'b01100000;
font_rom[1556] <= 8'b00001100;
font_rom[1557] <= 8'b11000000;
font_rom[1558] <= 8'b00001100;
font_rom[1559] <= 8'b11000000;
font_rom[1560] <= 8'b00000111;
font_rom[1561] <= 8'b11000000;
font_rom[1562] <= 8'b00000000;
font_rom[1563] <= 8'b00000000;
font_rom[1564] <= 8'b00000000;
font_rom[1565] <= 8'b00000000;
font_rom[1566] <= 8'b00000000;
font_rom[1567] <= 8'b00000000;
//ASCII 0x31 '1'
font_rom[1568] <= 8'b00000000;
font_rom[1569] <= 8'b00000000;
font_rom[1570] <= 8'b00000000;
font_rom[1571] <= 8'b00000000;
font_rom[1572] <= 8'b00000000;
font_rom[1573] <= 8'b00000000;
font_rom[1574] <= 8'b00000000;
font_rom[1575] <= 8'b00000000;
font_rom[1576] <= 8'b00000000;
font_rom[1577] <= 8'b00000000;
font_rom[1578] <= 8'b00000001;
font_rom[1579] <= 8'b10000000;
font_rom[1580] <= 8'b00000011;
font_rom[1581] <= 8'b10000000;
font_rom[1582] <= 8'b00000000;
font_rom[1583] <= 8'b10000000;
font_rom[1584] <= 8'b00000001;
font_rom[1585] <= 8'b10000000;
font_rom[1586] <= 8'b00000001;
font_rom[1587] <= 8'b10000000;
font_rom[1588] <= 8'b00000001;
font_rom[1589] <= 8'b10000000;
font_rom[1590] <= 8'b00000001;
font_rom[1591] <= 8'b10000000;
font_rom[1592] <= 8'b00000011;
font_rom[1593] <= 8'b11000000;
font_rom[1594] <= 8'b00000000;
font_rom[1595] <= 8'b00000000;
font_rom[1596] <= 8'b00000000;
font_rom[1597] <= 8'b00000000;
font_rom[1598] <= 8'b00000000;
font_rom[1599] <= 8'b00000000;
//ASCII 0x32 '2'
font_rom[1600] <= 8'b00000000;
font_rom[1601] <= 8'b00000000;
font_rom[1602] <= 8'b00000000;
font_rom[1603] <= 8'b00000000;
font_rom[1604] <= 8'b00000000;
font_rom[1605] <= 8'b00000000;
font_rom[1606] <= 8'b00000000;
font_rom[1607] <= 8'b00000000;
font_rom[1608] <= 8'b00000000;
font_rom[1609] <= 8'b00000000;
font_rom[1610] <= 8'b00000111;
font_rom[1611] <= 8'b10000000;
font_rom[1612] <= 8'b00001100;
font_rom[1613] <= 8'b11000000;
font_rom[1614] <= 8'b00000000;
font_rom[1615] <= 8'b11000000;
font_rom[1616] <= 8'b00000001;
font_rom[1617] <= 8'b11000000;
font_rom[1618] <= 8'b00000011;
font_rom[1619] <= 8'b00000000;
font_rom[1620] <= 8'b00000110;
font_rom[1621] <= 8'b00000000;
font_rom[1622] <= 8'b00001100;
font_rom[1623] <= 8'b00000000;
font_rom[1624] <= 8'b00001111;
font_rom[1625] <= 8'b11000000;
font_rom[1626] <= 8'b00000000;
font_rom[1627] <= 8'b00000000;
font_rom[1628] <= 8'b00000000;
font_rom[1629] <= 8'b00000000;
font_rom[1630] <= 8'b00000000;
font_rom[1631] <= 8'b00000000;
//ASCII 0x33 '3'
font_rom[1632] <= 8'b00000000;
font_rom[1633] <= 8'b00000000;
font_rom[1634] <= 8'b00000000;
font_rom[1635] <= 8'b00000000;
font_rom[1636] <= 8'b00000000;
font_rom[1637] <= 8'b00000000;
font_rom[1638] <= 8'b00000000;
font_rom[1639] <= 8'b00000000;
font_rom[1640] <= 8'b00000000;
font_rom[1641] <= 8'b00000000;
font_rom[1642] <= 8'b00000111;
font_rom[1643] <= 8'b10000000;
font_rom[1644] <= 8'b00001100;
font_rom[1645] <= 8'b11000000;
font_rom[1646] <= 8'b00000000;
font_rom[1647] <= 8'b11000000;
font_rom[1648] <= 8'b00000011;
font_rom[1649] <= 8'b10000000;
font_rom[1650] <= 8'b00000000;
font_rom[1651] <= 8'b11000000;
font_rom[1652] <= 8'b00000000;
font_rom[1653] <= 8'b11000000;
font_rom[1654] <= 8'b00001100;
font_rom[1655] <= 8'b11000000;
font_rom[1656] <= 8'b00000111;
font_rom[1657] <= 8'b10000000;
font_rom[1658] <= 8'b00000000;
font_rom[1659] <= 8'b00000000;
font_rom[1660] <= 8'b00000000;
font_rom[1661] <= 8'b00000000;
font_rom[1662] <= 8'b00000000;
font_rom[1663] <= 8'b00000000;
//ASCII 0x34 '4'
font_rom[1664] <= 8'b00000000;
font_rom[1665] <= 8'b00000000;
font_rom[1666] <= 8'b00000000;
font_rom[1667] <= 8'b00000000;
font_rom[1668] <= 8'b00000000;
font_rom[1669] <= 8'b00000000;
font_rom[1670] <= 8'b00000000;
font_rom[1671] <= 8'b00000000;
font_rom[1672] <= 8'b00000000;
font_rom[1673] <= 8'b00000000;
font_rom[1674] <= 8'b00000001;
font_rom[1675] <= 8'b10000000;
font_rom[1676] <= 8'b00000011;
font_rom[1677] <= 8'b10000000;
font_rom[1678] <= 8'b00000011;
font_rom[1679] <= 8'b10000000;
font_rom[1680] <= 8'b00000110;
font_rom[1681] <= 8'b10000000;
font_rom[1682] <= 8'b00001100;
font_rom[1683] <= 8'b10000000;
font_rom[1684] <= 8'b00001111;
font_rom[1685] <= 8'b11100000;
font_rom[1686] <= 8'b00000000;
font_rom[1687] <= 8'b10000000;
font_rom[1688] <= 8'b00000000;
font_rom[1689] <= 8'b10000000;
font_rom[1690] <= 8'b00000000;
font_rom[1691] <= 8'b00000000;
font_rom[1692] <= 8'b00000000;
font_rom[1693] <= 8'b00000000;
font_rom[1694] <= 8'b00000000;
font_rom[1695] <= 8'b00000000;
//ASCII 0x35 '5'
font_rom[1696] <= 8'b00000000;
font_rom[1697] <= 8'b00000000;
font_rom[1698] <= 8'b00000000;
font_rom[1699] <= 8'b00000000;
font_rom[1700] <= 8'b00000000;
font_rom[1701] <= 8'b00000000;
font_rom[1702] <= 8'b00000000;
font_rom[1703] <= 8'b00000000;
font_rom[1704] <= 8'b00000000;
font_rom[1705] <= 8'b00000000;
font_rom[1706] <= 8'b00001111;
font_rom[1707] <= 8'b11000000;
font_rom[1708] <= 8'b00001100;
font_rom[1709] <= 8'b00000000;
font_rom[1710] <= 8'b00001111;
font_rom[1711] <= 8'b11000000;
font_rom[1712] <= 8'b00001100;
font_rom[1713] <= 8'b11000000;
font_rom[1714] <= 8'b00000000;
font_rom[1715] <= 8'b01100000;
font_rom[1716] <= 8'b00000000;
font_rom[1717] <= 8'b01100000;
font_rom[1718] <= 8'b00001100;
font_rom[1719] <= 8'b11000000;
font_rom[1720] <= 8'b00000111;
font_rom[1721] <= 8'b10000000;
font_rom[1722] <= 8'b00000000;
font_rom[1723] <= 8'b00000000;
font_rom[1724] <= 8'b00000000;
font_rom[1725] <= 8'b00000000;
font_rom[1726] <= 8'b00000000;
font_rom[1727] <= 8'b00000000;
//ASCII 0x36 '6'
font_rom[1728] <= 8'b00000000;
font_rom[1729] <= 8'b00000000;
font_rom[1730] <= 8'b00000000;
font_rom[1731] <= 8'b00000000;
font_rom[1732] <= 8'b00000000;
font_rom[1733] <= 8'b00000000;
font_rom[1734] <= 8'b00000000;
font_rom[1735] <= 8'b00000000;
font_rom[1736] <= 8'b00000000;
font_rom[1737] <= 8'b00000000;
font_rom[1738] <= 8'b00000011;
font_rom[1739] <= 8'b10000000;
font_rom[1740] <= 8'b00000111;
font_rom[1741] <= 8'b00000000;
font_rom[1742] <= 8'b00000110;
font_rom[1743] <= 8'b00000000;
font_rom[1744] <= 8'b00001111;
font_rom[1745] <= 8'b10000000;
font_rom[1746] <= 8'b00001100;
font_rom[1747] <= 8'b11000000;
font_rom[1748] <= 8'b00001100;
font_rom[1749] <= 8'b11000000;
font_rom[1750] <= 8'b00001100;
font_rom[1751] <= 8'b11000000;
font_rom[1752] <= 8'b00000111;
font_rom[1753] <= 8'b10000000;
font_rom[1754] <= 8'b00000000;
font_rom[1755] <= 8'b00000000;
font_rom[1756] <= 8'b00000000;
font_rom[1757] <= 8'b00000000;
font_rom[1758] <= 8'b00000000;
font_rom[1759] <= 8'b00000000;
//ASCII 0x37 '7'
font_rom[1760] <= 8'b00000000;
font_rom[1761] <= 8'b00000000;
font_rom[1762] <= 8'b00000000;
font_rom[1763] <= 8'b00000000;
font_rom[1764] <= 8'b00000000;
font_rom[1765] <= 8'b00000000;
font_rom[1766] <= 8'b00000000;
font_rom[1767] <= 8'b00000000;
font_rom[1768] <= 8'b00000000;
font_rom[1769] <= 8'b00000000;
font_rom[1770] <= 8'b00001111;
font_rom[1771] <= 8'b11100000;
font_rom[1772] <= 8'b00000000;
font_rom[1773] <= 8'b11000000;
font_rom[1774] <= 8'b00000001;
font_rom[1775] <= 8'b10000000;
font_rom[1776] <= 8'b00000011;
font_rom[1777] <= 8'b00000000;
font_rom[1778] <= 8'b00000011;
font_rom[1779] <= 8'b00000000;
font_rom[1780] <= 8'b00000011;
font_rom[1781] <= 8'b00000000;
font_rom[1782] <= 8'b00000110;
font_rom[1783] <= 8'b00000000;
font_rom[1784] <= 8'b00000110;
font_rom[1785] <= 8'b00000000;
font_rom[1786] <= 8'b00000000;
font_rom[1787] <= 8'b00000000;
font_rom[1788] <= 8'b00000000;
font_rom[1789] <= 8'b00000000;
font_rom[1790] <= 8'b00000000;
font_rom[1791] <= 8'b00000000;
//ASCII 0x38 '8'
font_rom[1792] <= 8'b00000000;
font_rom[1793] <= 8'b00000000;
font_rom[1794] <= 8'b00000000;
font_rom[1795] <= 8'b00000000;
font_rom[1796] <= 8'b00000000;
font_rom[1797] <= 8'b00000000;
font_rom[1798] <= 8'b00000000;
font_rom[1799] <= 8'b00000000;
font_rom[1800] <= 8'b00000000;
font_rom[1801] <= 8'b00000000;
font_rom[1802] <= 8'b00000111;
font_rom[1803] <= 8'b10000000;
font_rom[1804] <= 8'b00001100;
font_rom[1805] <= 8'b11000000;
font_rom[1806] <= 8'b00001100;
font_rom[1807] <= 8'b11000000;
font_rom[1808] <= 8'b00000111;
font_rom[1809] <= 8'b10000000;
font_rom[1810] <= 8'b00001100;
font_rom[1811] <= 8'b11000000;
font_rom[1812] <= 8'b00001100;
font_rom[1813] <= 8'b11000000;
font_rom[1814] <= 8'b00001100;
font_rom[1815] <= 8'b11000000;
font_rom[1816] <= 8'b00000111;
font_rom[1817] <= 8'b10000000;
font_rom[1818] <= 8'b00000000;
font_rom[1819] <= 8'b00000000;
font_rom[1820] <= 8'b00000000;
font_rom[1821] <= 8'b00000000;
font_rom[1822] <= 8'b00000000;
font_rom[1823] <= 8'b00000000;
//ASCII 0x39 '9'
font_rom[1824] <= 8'b00000000;
font_rom[1825] <= 8'b00000000;
font_rom[1826] <= 8'b00000000;
font_rom[1827] <= 8'b00000000;
font_rom[1828] <= 8'b00000000;
font_rom[1829] <= 8'b00000000;
font_rom[1830] <= 8'b00000000;
font_rom[1831] <= 8'b00000000;
font_rom[1832] <= 8'b00000000;
font_rom[1833] <= 8'b00000000;
font_rom[1834] <= 8'b00000111;
font_rom[1835] <= 8'b10000000;
font_rom[1836] <= 8'b00001100;
font_rom[1837] <= 8'b11000000;
font_rom[1838] <= 8'b00001100;
font_rom[1839] <= 8'b01100000;
font_rom[1840] <= 8'b00001100;
font_rom[1841] <= 8'b01100000;
font_rom[1842] <= 8'b00000111;
font_rom[1843] <= 8'b11000000;
font_rom[1844] <= 8'b00000000;
font_rom[1845] <= 8'b11000000;
font_rom[1846] <= 8'b00000011;
font_rom[1847] <= 8'b10000000;
font_rom[1848] <= 8'b00001110;
font_rom[1849] <= 8'b00000000;
font_rom[1850] <= 8'b00000000;
font_rom[1851] <= 8'b00000000;
font_rom[1852] <= 8'b00000000;
font_rom[1853] <= 8'b00000000;
font_rom[1854] <= 8'b00000000;
font_rom[1855] <= 8'b00000000;
//ASCII 0x3A ':'
font_rom[1856] <= 8'b00000000;
font_rom[1857] <= 8'b00000000;
font_rom[1858] <= 8'b00000000;
font_rom[1859] <= 8'b00000000;
font_rom[1860] <= 8'b00000000;
font_rom[1861] <= 8'b00000000;
font_rom[1862] <= 8'b00000000;
font_rom[1863] <= 8'b00000000;
font_rom[1864] <= 8'b00000000;
font_rom[1865] <= 8'b00000000;
font_rom[1866] <= 8'b00000000;
font_rom[1867] <= 8'b00000000;
font_rom[1868] <= 8'b00000000;
font_rom[1869] <= 8'b00000000;
font_rom[1870] <= 8'b00000011;
font_rom[1871] <= 8'b00000000;
font_rom[1872] <= 8'b00000000;
font_rom[1873] <= 8'b00000000;
font_rom[1874] <= 8'b00000000;
font_rom[1875] <= 8'b00000000;
font_rom[1876] <= 8'b00000000;
font_rom[1877] <= 8'b00000000;
font_rom[1878] <= 8'b00000011;
font_rom[1879] <= 8'b00000000;
font_rom[1880] <= 8'b00000000;
font_rom[1881] <= 8'b00000000;
font_rom[1882] <= 8'b00000000;
font_rom[1883] <= 8'b00000000;
font_rom[1884] <= 8'b00000000;
font_rom[1885] <= 8'b00000000;
font_rom[1886] <= 8'b00000000;
font_rom[1887] <= 8'b00000000;
//ASCII 0x3B ';'
font_rom[1888] <= 8'b00000000;
font_rom[1889] <= 8'b00000000;
font_rom[1890] <= 8'b00000000;
font_rom[1891] <= 8'b00000000;
font_rom[1892] <= 8'b00000000;
font_rom[1893] <= 8'b00000000;
font_rom[1894] <= 8'b00000000;
font_rom[1895] <= 8'b00000000;
font_rom[1896] <= 8'b00000000;
font_rom[1897] <= 8'b00000000;
font_rom[1898] <= 8'b00000000;
font_rom[1899] <= 8'b00000000;
font_rom[1900] <= 8'b00000000;
font_rom[1901] <= 8'b00000000;
font_rom[1902] <= 8'b00000011;
font_rom[1903] <= 8'b00000000;
font_rom[1904] <= 8'b00000000;
font_rom[1905] <= 8'b00000000;
font_rom[1906] <= 8'b00000000;
font_rom[1907] <= 8'b00000000;
font_rom[1908] <= 8'b00000000;
font_rom[1909] <= 8'b00000000;
font_rom[1910] <= 8'b00000000;
font_rom[1911] <= 8'b00000000;
font_rom[1912] <= 8'b00000011;
font_rom[1913] <= 8'b00000000;
font_rom[1914] <= 8'b00000010;
font_rom[1915] <= 8'b00000000;
font_rom[1916] <= 8'b00000000;
font_rom[1917] <= 8'b00000000;
font_rom[1918] <= 8'b00000000;
font_rom[1919] <= 8'b00000000;
//ASCII 0x3C '<'
font_rom[1920] <= 8'b00000000;
font_rom[1921] <= 8'b00000000;
font_rom[1922] <= 8'b00000000;
font_rom[1923] <= 8'b00000000;
font_rom[1924] <= 8'b00000000;
font_rom[1925] <= 8'b00000000;
font_rom[1926] <= 8'b00000000;
font_rom[1927] <= 8'b00000000;
font_rom[1928] <= 8'b00000000;
font_rom[1929] <= 8'b00000000;
font_rom[1930] <= 8'b00000000;
font_rom[1931] <= 8'b00000000;
font_rom[1932] <= 8'b00000000;
font_rom[1933] <= 8'b00000000;
font_rom[1934] <= 8'b00000001;
font_rom[1935] <= 8'b10000000;
font_rom[1936] <= 8'b00000011;
font_rom[1937] <= 8'b10000000;
font_rom[1938] <= 8'b00000111;
font_rom[1939] <= 8'b00000000;
font_rom[1940] <= 8'b00000011;
font_rom[1941] <= 8'b00000000;
font_rom[1942] <= 8'b00000001;
font_rom[1943] <= 8'b10000000;
font_rom[1944] <= 8'b00000000;
font_rom[1945] <= 8'b00000000;
font_rom[1946] <= 8'b00000000;
font_rom[1947] <= 8'b00000000;
font_rom[1948] <= 8'b00000000;
font_rom[1949] <= 8'b00000000;
font_rom[1950] <= 8'b00000000;
font_rom[1951] <= 8'b00000000;
//ASCII 0x3D '='
font_rom[1952] <= 8'b00000000;
font_rom[1953] <= 8'b00000000;
font_rom[1954] <= 8'b00000000;
font_rom[1955] <= 8'b00000000;
font_rom[1956] <= 8'b00000000;
font_rom[1957] <= 8'b00000000;
font_rom[1958] <= 8'b00000000;
font_rom[1959] <= 8'b00000000;
font_rom[1960] <= 8'b00000000;
font_rom[1961] <= 8'b00000000;
font_rom[1962] <= 8'b00000000;
font_rom[1963] <= 8'b00000000;
font_rom[1964] <= 8'b00000000;
font_rom[1965] <= 8'b00000000;
font_rom[1966] <= 8'b00000111;
font_rom[1967] <= 8'b11000000;
font_rom[1968] <= 8'b00000000;
font_rom[1969] <= 8'b00000000;
font_rom[1970] <= 8'b00000000;
font_rom[1971] <= 8'b00000000;
font_rom[1972] <= 8'b00000111;
font_rom[1973] <= 8'b11000000;
font_rom[1974] <= 8'b00000000;
font_rom[1975] <= 8'b00000000;
font_rom[1976] <= 8'b00000000;
font_rom[1977] <= 8'b00000000;
font_rom[1978] <= 8'b00000000;
font_rom[1979] <= 8'b00000000;
font_rom[1980] <= 8'b00000000;
font_rom[1981] <= 8'b00000000;
font_rom[1982] <= 8'b00000000;
font_rom[1983] <= 8'b00000000;
//ASCII 0x3E '>'
font_rom[1984] <= 8'b00000000;
font_rom[1985] <= 8'b00000000;
font_rom[1986] <= 8'b00000000;
font_rom[1987] <= 8'b00000000;
font_rom[1988] <= 8'b00000000;
font_rom[1989] <= 8'b00000000;
font_rom[1990] <= 8'b00000000;
font_rom[1991] <= 8'b00000000;
font_rom[1992] <= 8'b00000000;
font_rom[1993] <= 8'b00000000;
font_rom[1994] <= 8'b00000000;
font_rom[1995] <= 8'b00000000;
font_rom[1996] <= 8'b00000000;
font_rom[1997] <= 8'b00000000;
font_rom[1998] <= 8'b00000011;
font_rom[1999] <= 8'b00000000;
font_rom[2000] <= 8'b00000001;
font_rom[2001] <= 8'b10000000;
font_rom[2002] <= 8'b00000000;
font_rom[2003] <= 8'b11000000;
font_rom[2004] <= 8'b00000001;
font_rom[2005] <= 8'b10000000;
font_rom[2006] <= 8'b00000011;
font_rom[2007] <= 8'b00000000;
font_rom[2008] <= 8'b00000000;
font_rom[2009] <= 8'b00000000;
font_rom[2010] <= 8'b00000000;
font_rom[2011] <= 8'b00000000;
font_rom[2012] <= 8'b00000000;
font_rom[2013] <= 8'b00000000;
font_rom[2014] <= 8'b00000000;
font_rom[2015] <= 8'b00000000;
//ASCII 0x3F '?'
font_rom[2016] <= 8'b00000000;
font_rom[2017] <= 8'b00000000;
font_rom[2018] <= 8'b00000000;
font_rom[2019] <= 8'b00000000;
font_rom[2020] <= 8'b00000000;
font_rom[2021] <= 8'b00000000;
font_rom[2022] <= 8'b00000000;
font_rom[2023] <= 8'b00000000;
font_rom[2024] <= 8'b00000000;
font_rom[2025] <= 8'b00000000;
font_rom[2026] <= 8'b00000111;
font_rom[2027] <= 8'b10000000;
font_rom[2028] <= 8'b00000000;
font_rom[2029] <= 8'b11000000;
font_rom[2030] <= 8'b00000000;
font_rom[2031] <= 8'b01000000;
font_rom[2032] <= 8'b00000000;
font_rom[2033] <= 8'b11000000;
font_rom[2034] <= 8'b00000011;
font_rom[2035] <= 8'b10000000;
font_rom[2036] <= 8'b00000011;
font_rom[2037] <= 8'b00000000;
font_rom[2038] <= 8'b00000000;
font_rom[2039] <= 8'b00000000;
font_rom[2040] <= 8'b00000110;
font_rom[2041] <= 8'b00000000;
font_rom[2042] <= 8'b00000000;
font_rom[2043] <= 8'b00000000;
font_rom[2044] <= 8'b00000000;
font_rom[2045] <= 8'b00000000;
font_rom[2046] <= 8'b00000000;
font_rom[2047] <= 8'b00000000;
//ASCII 0x40 '@'
font_rom[2048] <= 8'b00000000;
font_rom[2049] <= 8'b00000000;
font_rom[2050] <= 8'b00000000;
font_rom[2051] <= 8'b00000000;
font_rom[2052] <= 8'b00000000;
font_rom[2053] <= 8'b00000000;
font_rom[2054] <= 8'b00000000;
font_rom[2055] <= 8'b00000000;
font_rom[2056] <= 8'b00000111;
font_rom[2057] <= 8'b11000000;
font_rom[2058] <= 8'b00001100;
font_rom[2059] <= 8'b01100000;
font_rom[2060] <= 8'b00011011;
font_rom[2061] <= 8'b10110000;
font_rom[2062] <= 8'b00011111;
font_rom[2063] <= 8'b10110000;
font_rom[2064] <= 8'b00011111;
font_rom[2065] <= 8'b10110000;
font_rom[2066] <= 8'b00011111;
font_rom[2067] <= 8'b11110000;
font_rom[2068] <= 8'b00011000;
font_rom[2069] <= 8'b00000000;
font_rom[2070] <= 8'b00001100;
font_rom[2071] <= 8'b01100000;
font_rom[2072] <= 8'b00000111;
font_rom[2073] <= 8'b11000000;
font_rom[2074] <= 8'b00000000;
font_rom[2075] <= 8'b00000000;
font_rom[2076] <= 8'b00000000;
font_rom[2077] <= 8'b00000000;
font_rom[2078] <= 8'b00000000;
font_rom[2079] <= 8'b00000000;
//ASCII 0x41 'A'
font_rom[2080] <= 8'b00000000;
font_rom[2081] <= 8'b00000000;
font_rom[2082] <= 8'b00000000;
font_rom[2083] <= 8'b00000000;
font_rom[2084] <= 8'b00000000;
font_rom[2085] <= 8'b00000000;
font_rom[2086] <= 8'b00000000;
font_rom[2087] <= 8'b00000000;
font_rom[2088] <= 8'b00000000;
font_rom[2089] <= 8'b00000000;
font_rom[2090] <= 8'b00000000;
font_rom[2091] <= 8'b11000000;
font_rom[2092] <= 8'b00000001;
font_rom[2093] <= 8'b11000000;
font_rom[2094] <= 8'b00000011;
font_rom[2095] <= 8'b11000000;
font_rom[2096] <= 8'b00000011;
font_rom[2097] <= 8'b11000000;
font_rom[2098] <= 8'b00000111;
font_rom[2099] <= 8'b11100000;
font_rom[2100] <= 8'b00000110;
font_rom[2101] <= 8'b01100000;
font_rom[2102] <= 8'b00001100;
font_rom[2103] <= 8'b01100000;
font_rom[2104] <= 8'b00001100;
font_rom[2105] <= 8'b01100000;
font_rom[2106] <= 8'b00000000;
font_rom[2107] <= 8'b00000000;
font_rom[2108] <= 8'b00000000;
font_rom[2109] <= 8'b00000000;
font_rom[2110] <= 8'b00000000;
font_rom[2111] <= 8'b00000000;
//ASCII 0x42 'B'
font_rom[2112] <= 8'b00000000;
font_rom[2113] <= 8'b00000000;
font_rom[2114] <= 8'b00000000;
font_rom[2115] <= 8'b00000000;
font_rom[2116] <= 8'b00000000;
font_rom[2117] <= 8'b00000000;
font_rom[2118] <= 8'b00000000;
font_rom[2119] <= 8'b00000000;
font_rom[2120] <= 8'b00000000;
font_rom[2121] <= 8'b00000000;
font_rom[2122] <= 8'b00000111;
font_rom[2123] <= 8'b10000000;
font_rom[2124] <= 8'b00001100;
font_rom[2125] <= 8'b11000000;
font_rom[2126] <= 8'b00001100;
font_rom[2127] <= 8'b11000000;
font_rom[2128] <= 8'b00001100;
font_rom[2129] <= 8'b11000000;
font_rom[2130] <= 8'b00001111;
font_rom[2131] <= 8'b10000000;
font_rom[2132] <= 8'b00001100;
font_rom[2133] <= 8'b11100000;
font_rom[2134] <= 8'b00001100;
font_rom[2135] <= 8'b11000000;
font_rom[2136] <= 8'b00001111;
font_rom[2137] <= 8'b10000000;
font_rom[2138] <= 8'b00000000;
font_rom[2139] <= 8'b00000000;
font_rom[2140] <= 8'b00000000;
font_rom[2141] <= 8'b00000000;
font_rom[2142] <= 8'b00000000;
font_rom[2143] <= 8'b00000000;
//ASCII 0x43 'C'
font_rom[2144] <= 8'b00000000;
font_rom[2145] <= 8'b00000000;
font_rom[2146] <= 8'b00000000;
font_rom[2147] <= 8'b00000000;
font_rom[2148] <= 8'b00000000;
font_rom[2149] <= 8'b00000000;
font_rom[2150] <= 8'b00000000;
font_rom[2151] <= 8'b00000000;
font_rom[2152] <= 8'b00000000;
font_rom[2153] <= 8'b00000000;
font_rom[2154] <= 8'b00000011;
font_rom[2155] <= 8'b11100000;
font_rom[2156] <= 8'b00000111;
font_rom[2157] <= 8'b01100000;
font_rom[2158] <= 8'b00000110;
font_rom[2159] <= 8'b00000000;
font_rom[2160] <= 8'b00001100;
font_rom[2161] <= 8'b00000000;
font_rom[2162] <= 8'b00001100;
font_rom[2163] <= 8'b00000000;
font_rom[2164] <= 8'b00001100;
font_rom[2165] <= 8'b00000000;
font_rom[2166] <= 8'b00001100;
font_rom[2167] <= 8'b11000000;
font_rom[2168] <= 8'b00000111;
font_rom[2169] <= 8'b10000000;
font_rom[2170] <= 8'b00000000;
font_rom[2171] <= 8'b00000000;
font_rom[2172] <= 8'b00000000;
font_rom[2173] <= 8'b00000000;
font_rom[2174] <= 8'b00000000;
font_rom[2175] <= 8'b00000000;
//ASCII 0x44 'D'
font_rom[2176] <= 8'b00000000;
font_rom[2177] <= 8'b00000000;
font_rom[2178] <= 8'b00000000;
font_rom[2179] <= 8'b00000000;
font_rom[2180] <= 8'b00000000;
font_rom[2181] <= 8'b00000000;
font_rom[2182] <= 8'b00000000;
font_rom[2183] <= 8'b00000000;
font_rom[2184] <= 8'b00000000;
font_rom[2185] <= 8'b00000000;
font_rom[2186] <= 8'b00001110;
font_rom[2187] <= 8'b00000000;
font_rom[2188] <= 8'b00001111;
font_rom[2189] <= 8'b10000000;
font_rom[2190] <= 8'b00001100;
font_rom[2191] <= 8'b11100000;
font_rom[2192] <= 8'b00001100;
font_rom[2193] <= 8'b01100000;
font_rom[2194] <= 8'b00001100;
font_rom[2195] <= 8'b00100000;
font_rom[2196] <= 8'b00001100;
font_rom[2197] <= 8'b01100000;
font_rom[2198] <= 8'b00001100;
font_rom[2199] <= 8'b01100000;
font_rom[2200] <= 8'b00000111;
font_rom[2201] <= 8'b11000000;
font_rom[2202] <= 8'b00000000;
font_rom[2203] <= 8'b00000000;
font_rom[2204] <= 8'b00000000;
font_rom[2205] <= 8'b00000000;
font_rom[2206] <= 8'b00000000;
font_rom[2207] <= 8'b00000000;
//ASCII 0x45 'E'
font_rom[2208] <= 8'b00000000;
font_rom[2209] <= 8'b00000000;
font_rom[2210] <= 8'b00000000;
font_rom[2211] <= 8'b00000000;
font_rom[2212] <= 8'b00000000;
font_rom[2213] <= 8'b00000000;
font_rom[2214] <= 8'b00000000;
font_rom[2215] <= 8'b00000000;
font_rom[2216] <= 8'b00000000;
font_rom[2217] <= 8'b00000000;
font_rom[2218] <= 8'b00001111;
font_rom[2219] <= 8'b11100000;
font_rom[2220] <= 8'b00001100;
font_rom[2221] <= 8'b00000000;
font_rom[2222] <= 8'b00001100;
font_rom[2223] <= 8'b00000000;
font_rom[2224] <= 8'b00001111;
font_rom[2225] <= 8'b11000000;
font_rom[2226] <= 8'b00001100;
font_rom[2227] <= 8'b00000000;
font_rom[2228] <= 8'b00001100;
font_rom[2229] <= 8'b00000000;
font_rom[2230] <= 8'b00001100;
font_rom[2231] <= 8'b00000000;
font_rom[2232] <= 8'b00001111;
font_rom[2233] <= 8'b11000000;
font_rom[2234] <= 8'b00000000;
font_rom[2235] <= 8'b00000000;
font_rom[2236] <= 8'b00000000;
font_rom[2237] <= 8'b00000000;
font_rom[2238] <= 8'b00000000;
font_rom[2239] <= 8'b00000000;
//ASCII 0x46 'F'
font_rom[2240] <= 8'b00000000;
font_rom[2241] <= 8'b00000000;
font_rom[2242] <= 8'b00000000;
font_rom[2243] <= 8'b00000000;
font_rom[2244] <= 8'b00000000;
font_rom[2245] <= 8'b00000000;
font_rom[2246] <= 8'b00000000;
font_rom[2247] <= 8'b00000000;
font_rom[2248] <= 8'b00000000;
font_rom[2249] <= 8'b00000000;
font_rom[2250] <= 8'b00000111;
font_rom[2251] <= 8'b11100000;
font_rom[2252] <= 8'b00000110;
font_rom[2253] <= 8'b00000000;
font_rom[2254] <= 8'b00000110;
font_rom[2255] <= 8'b00000000;
font_rom[2256] <= 8'b00000111;
font_rom[2257] <= 8'b11100000;
font_rom[2258] <= 8'b00000110;
font_rom[2259] <= 8'b00000000;
font_rom[2260] <= 8'b00000110;
font_rom[2261] <= 8'b00000000;
font_rom[2262] <= 8'b00000110;
font_rom[2263] <= 8'b00000000;
font_rom[2264] <= 8'b00000110;
font_rom[2265] <= 8'b00000000;
font_rom[2266] <= 8'b00000000;
font_rom[2267] <= 8'b00000000;
font_rom[2268] <= 8'b00000000;
font_rom[2269] <= 8'b00000000;
font_rom[2270] <= 8'b00000000;
font_rom[2271] <= 8'b00000000;
//ASCII 0x47 'G'
font_rom[2272] <= 8'b00000000;
font_rom[2273] <= 8'b00000000;
font_rom[2274] <= 8'b00000000;
font_rom[2275] <= 8'b00000000;
font_rom[2276] <= 8'b00000000;
font_rom[2277] <= 8'b00000000;
font_rom[2278] <= 8'b00000000;
font_rom[2279] <= 8'b00000000;
font_rom[2280] <= 8'b00000000;
font_rom[2281] <= 8'b00000000;
font_rom[2282] <= 8'b00000011;
font_rom[2283] <= 8'b11000000;
font_rom[2284] <= 8'b00000110;
font_rom[2285] <= 8'b01100000;
font_rom[2286] <= 8'b00000110;
font_rom[2287] <= 8'b00000000;
font_rom[2288] <= 8'b00001100;
font_rom[2289] <= 8'b00000000;
font_rom[2290] <= 8'b00001111;
font_rom[2291] <= 8'b11100000;
font_rom[2292] <= 8'b00001100;
font_rom[2293] <= 8'b01100000;
font_rom[2294] <= 8'b00001100;
font_rom[2295] <= 8'b01100000;
font_rom[2296] <= 8'b00000111;
font_rom[2297] <= 8'b11000000;
font_rom[2298] <= 8'b00000000;
font_rom[2299] <= 8'b00000000;
font_rom[2300] <= 8'b00000000;
font_rom[2301] <= 8'b00000000;
font_rom[2302] <= 8'b00000000;
font_rom[2303] <= 8'b00000000;
//ASCII 0x48 'H'
font_rom[2304] <= 8'b00000000;
font_rom[2305] <= 8'b00000000;
font_rom[2306] <= 8'b00000000;
font_rom[2307] <= 8'b00000000;
font_rom[2308] <= 8'b00000000;
font_rom[2309] <= 8'b00000000;
font_rom[2310] <= 8'b00000000;
font_rom[2311] <= 8'b00000000;
font_rom[2312] <= 8'b00000000;
font_rom[2313] <= 8'b00000000;
font_rom[2314] <= 8'b00001100;
font_rom[2315] <= 8'b00110000;
font_rom[2316] <= 8'b00001100;
font_rom[2317] <= 8'b00100000;
font_rom[2318] <= 8'b00001100;
font_rom[2319] <= 8'b00100000;
font_rom[2320] <= 8'b00001111;
font_rom[2321] <= 8'b11100000;
font_rom[2322] <= 8'b00001110;
font_rom[2323] <= 8'b01100000;
font_rom[2324] <= 8'b00001100;
font_rom[2325] <= 8'b01100000;
font_rom[2326] <= 8'b00001100;
font_rom[2327] <= 8'b01100000;
font_rom[2328] <= 8'b00001100;
font_rom[2329] <= 8'b01100000;
font_rom[2330] <= 8'b00000000;
font_rom[2331] <= 8'b00000000;
font_rom[2332] <= 8'b00000000;
font_rom[2333] <= 8'b00000000;
font_rom[2334] <= 8'b00000000;
font_rom[2335] <= 8'b00000000;
//ASCII 0x49 'I'
font_rom[2336] <= 8'b00000000;
font_rom[2337] <= 8'b00000000;
font_rom[2338] <= 8'b00000000;
font_rom[2339] <= 8'b00000000;
font_rom[2340] <= 8'b00000000;
font_rom[2341] <= 8'b00000000;
font_rom[2342] <= 8'b00000000;
font_rom[2343] <= 8'b00000000;
font_rom[2344] <= 8'b00000000;
font_rom[2345] <= 8'b00000000;
font_rom[2346] <= 8'b00000111;
font_rom[2347] <= 8'b11100000;
font_rom[2348] <= 8'b00000001;
font_rom[2349] <= 8'b00000000;
font_rom[2350] <= 8'b00000011;
font_rom[2351] <= 8'b00000000;
font_rom[2352] <= 8'b00000011;
font_rom[2353] <= 8'b00000000;
font_rom[2354] <= 8'b00000011;
font_rom[2355] <= 8'b00000000;
font_rom[2356] <= 8'b00000001;
font_rom[2357] <= 8'b00000000;
font_rom[2358] <= 8'b00000001;
font_rom[2359] <= 8'b00000000;
font_rom[2360] <= 8'b00000111;
font_rom[2361] <= 8'b11000000;
font_rom[2362] <= 8'b00000000;
font_rom[2363] <= 8'b00000000;
font_rom[2364] <= 8'b00000000;
font_rom[2365] <= 8'b00000000;
font_rom[2366] <= 8'b00000000;
font_rom[2367] <= 8'b00000000;
//ASCII 0x4A 'J'
font_rom[2368] <= 8'b00000000;
font_rom[2369] <= 8'b00000000;
font_rom[2370] <= 8'b00000000;
font_rom[2371] <= 8'b00000000;
font_rom[2372] <= 8'b00000000;
font_rom[2373] <= 8'b00000000;
font_rom[2374] <= 8'b00000000;
font_rom[2375] <= 8'b00000000;
font_rom[2376] <= 8'b00000000;
font_rom[2377] <= 8'b00000000;
font_rom[2378] <= 8'b00000111;
font_rom[2379] <= 8'b11100000;
font_rom[2380] <= 8'b00000001;
font_rom[2381] <= 8'b10000000;
font_rom[2382] <= 8'b00000001;
font_rom[2383] <= 8'b10000000;
font_rom[2384] <= 8'b00000001;
font_rom[2385] <= 8'b10000000;
font_rom[2386] <= 8'b00000001;
font_rom[2387] <= 8'b10000000;
font_rom[2388] <= 8'b00001101;
font_rom[2389] <= 8'b10000000;
font_rom[2390] <= 8'b00001101;
font_rom[2391] <= 8'b10000000;
font_rom[2392] <= 8'b00000111;
font_rom[2393] <= 8'b00000000;
font_rom[2394] <= 8'b00000000;
font_rom[2395] <= 8'b00000000;
font_rom[2396] <= 8'b00000000;
font_rom[2397] <= 8'b00000000;
font_rom[2398] <= 8'b00000000;
font_rom[2399] <= 8'b00000000;
//ASCII 0x4B 'K'
font_rom[2400] <= 8'b00000000;
font_rom[2401] <= 8'b00000000;
font_rom[2402] <= 8'b00000000;
font_rom[2403] <= 8'b00000000;
font_rom[2404] <= 8'b00000000;
font_rom[2405] <= 8'b00000000;
font_rom[2406] <= 8'b00000000;
font_rom[2407] <= 8'b00000000;
font_rom[2408] <= 8'b00000000;
font_rom[2409] <= 8'b00000000;
font_rom[2410] <= 8'b00000100;
font_rom[2411] <= 8'b11100000;
font_rom[2412] <= 8'b00000100;
font_rom[2413] <= 8'b11000000;
font_rom[2414] <= 8'b00000101;
font_rom[2415] <= 8'b10000000;
font_rom[2416] <= 8'b00000111;
font_rom[2417] <= 8'b00000000;
font_rom[2418] <= 8'b00000111;
font_rom[2419] <= 8'b00000000;
font_rom[2420] <= 8'b00000111;
font_rom[2421] <= 8'b10000000;
font_rom[2422] <= 8'b00000101;
font_rom[2423] <= 8'b11000000;
font_rom[2424] <= 8'b00000100;
font_rom[2425] <= 8'b11100000;
font_rom[2426] <= 8'b00000000;
font_rom[2427] <= 8'b00000000;
font_rom[2428] <= 8'b00000000;
font_rom[2429] <= 8'b00000000;
font_rom[2430] <= 8'b00000000;
font_rom[2431] <= 8'b00000000;
//ASCII 0x4C 'L'
font_rom[2432] <= 8'b00000000;
font_rom[2433] <= 8'b00000000;
font_rom[2434] <= 8'b00000000;
font_rom[2435] <= 8'b00000000;
font_rom[2436] <= 8'b00000000;
font_rom[2437] <= 8'b00000000;
font_rom[2438] <= 8'b00000000;
font_rom[2439] <= 8'b00000000;
font_rom[2440] <= 8'b00000000;
font_rom[2441] <= 8'b00000000;
font_rom[2442] <= 8'b00000110;
font_rom[2443] <= 8'b00000000;
font_rom[2444] <= 8'b00000110;
font_rom[2445] <= 8'b00000000;
font_rom[2446] <= 8'b00000110;
font_rom[2447] <= 8'b00000000;
font_rom[2448] <= 8'b00000110;
font_rom[2449] <= 8'b00000000;
font_rom[2450] <= 8'b00000110;
font_rom[2451] <= 8'b00000000;
font_rom[2452] <= 8'b00000110;
font_rom[2453] <= 8'b00000000;
font_rom[2454] <= 8'b00000110;
font_rom[2455] <= 8'b00000000;
font_rom[2456] <= 8'b00000111;
font_rom[2457] <= 8'b11100000;
font_rom[2458] <= 8'b00000000;
font_rom[2459] <= 8'b00000000;
font_rom[2460] <= 8'b00000000;
font_rom[2461] <= 8'b00000000;
font_rom[2462] <= 8'b00000000;
font_rom[2463] <= 8'b00000000;
//ASCII 0x4D 'M'
font_rom[2464] <= 8'b00000000;
font_rom[2465] <= 8'b00000000;
font_rom[2466] <= 8'b00000000;
font_rom[2467] <= 8'b00000000;
font_rom[2468] <= 8'b00000000;
font_rom[2469] <= 8'b00000000;
font_rom[2470] <= 8'b00000000;
font_rom[2471] <= 8'b00000000;
font_rom[2472] <= 8'b00000000;
font_rom[2473] <= 8'b00000000;
font_rom[2474] <= 8'b00000110;
font_rom[2475] <= 8'b01100000;
font_rom[2476] <= 8'b00001110;
font_rom[2477] <= 8'b01100000;
font_rom[2478] <= 8'b00001110;
font_rom[2479] <= 8'b11100000;
font_rom[2480] <= 8'b00001110;
font_rom[2481] <= 8'b11100000;
font_rom[2482] <= 8'b00001110;
font_rom[2483] <= 8'b11110000;
font_rom[2484] <= 8'b00011011;
font_rom[2485] <= 8'b10110000;
font_rom[2486] <= 8'b00011011;
font_rom[2487] <= 8'b10110000;
font_rom[2488] <= 8'b00011011;
font_rom[2489] <= 8'b10110000;
font_rom[2490] <= 8'b00000000;
font_rom[2491] <= 8'b00000000;
font_rom[2492] <= 8'b00000000;
font_rom[2493] <= 8'b00000000;
font_rom[2494] <= 8'b00000000;
font_rom[2495] <= 8'b00000000;
//ASCII 0x4E 'N'
font_rom[2496] <= 8'b00000000;
font_rom[2497] <= 8'b00000000;
font_rom[2498] <= 8'b00000000;
font_rom[2499] <= 8'b00000000;
font_rom[2500] <= 8'b00000000;
font_rom[2501] <= 8'b00000000;
font_rom[2502] <= 8'b00000000;
font_rom[2503] <= 8'b00000000;
font_rom[2504] <= 8'b00000000;
font_rom[2505] <= 8'b00000000;
font_rom[2506] <= 8'b00001100;
font_rom[2507] <= 8'b00110000;
font_rom[2508] <= 8'b00001110;
font_rom[2509] <= 8'b00110000;
font_rom[2510] <= 8'b00001111;
font_rom[2511] <= 8'b00011000;
font_rom[2512] <= 8'b00001111;
font_rom[2513] <= 8'b00011000;
font_rom[2514] <= 8'b00001101;
font_rom[2515] <= 8'b10011000;
font_rom[2516] <= 8'b00001100;
font_rom[2517] <= 8'b11011000;
font_rom[2518] <= 8'b00001100;
font_rom[2519] <= 8'b01111000;
font_rom[2520] <= 8'b00001100;
font_rom[2521] <= 8'b00110000;
font_rom[2522] <= 8'b00000000;
font_rom[2523] <= 8'b00000000;
font_rom[2524] <= 8'b00000000;
font_rom[2525] <= 8'b00000000;
font_rom[2526] <= 8'b00000000;
font_rom[2527] <= 8'b00000000;
//ASCII 0x4F 'O'
font_rom[2528] <= 8'b00000000;
font_rom[2529] <= 8'b00000000;
font_rom[2530] <= 8'b00000000;
font_rom[2531] <= 8'b00000000;
font_rom[2532] <= 8'b00000000;
font_rom[2533] <= 8'b00000000;
font_rom[2534] <= 8'b00000000;
font_rom[2535] <= 8'b00000000;
font_rom[2536] <= 8'b00000000;
font_rom[2537] <= 8'b00000000;
font_rom[2538] <= 8'b00000011;
font_rom[2539] <= 8'b11100000;
font_rom[2540] <= 8'b00000110;
font_rom[2541] <= 8'b00110000;
font_rom[2542] <= 8'b00001100;
font_rom[2543] <= 8'b00011000;
font_rom[2544] <= 8'b00001100;
font_rom[2545] <= 8'b00011000;
font_rom[2546] <= 8'b00001100;
font_rom[2547] <= 8'b00010000;
font_rom[2548] <= 8'b00001100;
font_rom[2549] <= 8'b00110000;
font_rom[2550] <= 8'b00001110;
font_rom[2551] <= 8'b01100000;
font_rom[2552] <= 8'b00000011;
font_rom[2553] <= 8'b11000000;
font_rom[2554] <= 8'b00000000;
font_rom[2555] <= 8'b00000000;
font_rom[2556] <= 8'b00000000;
font_rom[2557] <= 8'b00000000;
font_rom[2558] <= 8'b00000000;
font_rom[2559] <= 8'b00000000;
//ASCII 0x50 'P'
font_rom[2560] <= 8'b00000000;
font_rom[2561] <= 8'b00000000;
font_rom[2562] <= 8'b00000000;
font_rom[2563] <= 8'b00000000;
font_rom[2564] <= 8'b00000000;
font_rom[2565] <= 8'b00000000;
font_rom[2566] <= 8'b00000000;
font_rom[2567] <= 8'b00000000;
font_rom[2568] <= 8'b00000000;
font_rom[2569] <= 8'b00000000;
font_rom[2570] <= 8'b00000111;
font_rom[2571] <= 8'b10000000;
font_rom[2572] <= 8'b00000110;
font_rom[2573] <= 8'b11000000;
font_rom[2574] <= 8'b00000110;
font_rom[2575] <= 8'b01100000;
font_rom[2576] <= 8'b00000110;
font_rom[2577] <= 8'b01100000;
font_rom[2578] <= 8'b00000110;
font_rom[2579] <= 8'b11000000;
font_rom[2580] <= 8'b00000111;
font_rom[2581] <= 8'b10000000;
font_rom[2582] <= 8'b00000110;
font_rom[2583] <= 8'b00000000;
font_rom[2584] <= 8'b00000110;
font_rom[2585] <= 8'b00000000;
font_rom[2586] <= 8'b00000000;
font_rom[2587] <= 8'b00000000;
font_rom[2588] <= 8'b00000000;
font_rom[2589] <= 8'b00000000;
font_rom[2590] <= 8'b00000000;
font_rom[2591] <= 8'b00000000;
//ASCII 0x51 'Q'
font_rom[2592] <= 8'b00000000;
font_rom[2593] <= 8'b00000000;
font_rom[2594] <= 8'b00000000;
font_rom[2595] <= 8'b00000000;
font_rom[2596] <= 8'b00000000;
font_rom[2597] <= 8'b00000000;
font_rom[2598] <= 8'b00000000;
font_rom[2599] <= 8'b00000000;
font_rom[2600] <= 8'b00000000;
font_rom[2601] <= 8'b00000000;
font_rom[2602] <= 8'b00000111;
font_rom[2603] <= 8'b11100000;
font_rom[2604] <= 8'b00001100;
font_rom[2605] <= 8'b01110000;
font_rom[2606] <= 8'b00011000;
font_rom[2607] <= 8'b00110000;
font_rom[2608] <= 8'b00011000;
font_rom[2609] <= 8'b00010000;
font_rom[2610] <= 8'b00011000;
font_rom[2611] <= 8'b00011000;
font_rom[2612] <= 8'b00011001;
font_rom[2613] <= 8'b10110000;
font_rom[2614] <= 8'b00001101;
font_rom[2615] <= 8'b11110000;
font_rom[2616] <= 8'b00000111;
font_rom[2617] <= 8'b11100000;
font_rom[2618] <= 8'b00000000;
font_rom[2619] <= 8'b00110000;
font_rom[2620] <= 8'b00000000;
font_rom[2621] <= 8'b00011000;
font_rom[2622] <= 8'b00000000;
font_rom[2623] <= 8'b00000000;
//ASCII 0x52 'R'
font_rom[2624] <= 8'b00000000;
font_rom[2625] <= 8'b00000000;
font_rom[2626] <= 8'b00000000;
font_rom[2627] <= 8'b00000000;
font_rom[2628] <= 8'b00000000;
font_rom[2629] <= 8'b00000000;
font_rom[2630] <= 8'b00000000;
font_rom[2631] <= 8'b00000000;
font_rom[2632] <= 8'b00000000;
font_rom[2633] <= 8'b00000000;
font_rom[2634] <= 8'b00001111;
font_rom[2635] <= 8'b00000000;
font_rom[2636] <= 8'b00001101;
font_rom[2637] <= 8'b11000000;
font_rom[2638] <= 8'b00001100;
font_rom[2639] <= 8'b11000000;
font_rom[2640] <= 8'b00001100;
font_rom[2641] <= 8'b11000000;
font_rom[2642] <= 8'b00001111;
font_rom[2643] <= 8'b10000000;
font_rom[2644] <= 8'b00001111;
font_rom[2645] <= 8'b10000000;
font_rom[2646] <= 8'b00001100;
font_rom[2647] <= 8'b11000000;
font_rom[2648] <= 8'b00001100;
font_rom[2649] <= 8'b01100000;
font_rom[2650] <= 8'b00000000;
font_rom[2651] <= 8'b00000000;
font_rom[2652] <= 8'b00000000;
font_rom[2653] <= 8'b00000000;
font_rom[2654] <= 8'b00000000;
font_rom[2655] <= 8'b00000000;
//ASCII 0x53 'S'
font_rom[2656] <= 8'b00000000;
font_rom[2657] <= 8'b00000000;
font_rom[2658] <= 8'b00000000;
font_rom[2659] <= 8'b00000000;
font_rom[2660] <= 8'b00000000;
font_rom[2661] <= 8'b00000000;
font_rom[2662] <= 8'b00000000;
font_rom[2663] <= 8'b00000000;
font_rom[2664] <= 8'b00000000;
font_rom[2665] <= 8'b00000000;
font_rom[2666] <= 8'b00000011;
font_rom[2667] <= 8'b11100000;
font_rom[2668] <= 8'b00000110;
font_rom[2669] <= 8'b00000000;
font_rom[2670] <= 8'b00000110;
font_rom[2671] <= 8'b00000000;
font_rom[2672] <= 8'b00000111;
font_rom[2673] <= 8'b11000000;
font_rom[2674] <= 8'b00000000;
font_rom[2675] <= 8'b01100000;
font_rom[2676] <= 8'b00000000;
font_rom[2677] <= 8'b00100000;
font_rom[2678] <= 8'b00001100;
font_rom[2679] <= 8'b01100000;
font_rom[2680] <= 8'b00000111;
font_rom[2681] <= 8'b11000000;
font_rom[2682] <= 8'b00000000;
font_rom[2683] <= 8'b00000000;
font_rom[2684] <= 8'b00000000;
font_rom[2685] <= 8'b00000000;
font_rom[2686] <= 8'b00000000;
font_rom[2687] <= 8'b00000000;
//ASCII 0x54 'T'
font_rom[2688] <= 8'b00000000;
font_rom[2689] <= 8'b00000000;
font_rom[2690] <= 8'b00000000;
font_rom[2691] <= 8'b00000000;
font_rom[2692] <= 8'b00000000;
font_rom[2693] <= 8'b00000000;
font_rom[2694] <= 8'b00000000;
font_rom[2695] <= 8'b00000000;
font_rom[2696] <= 8'b00000000;
font_rom[2697] <= 8'b00000000;
font_rom[2698] <= 8'b00001111;
font_rom[2699] <= 8'b11110000;
font_rom[2700] <= 8'b00000011;
font_rom[2701] <= 8'b00000000;
font_rom[2702] <= 8'b00000011;
font_rom[2703] <= 8'b00000000;
font_rom[2704] <= 8'b00000001;
font_rom[2705] <= 8'b00000000;
font_rom[2706] <= 8'b00000001;
font_rom[2707] <= 8'b00000000;
font_rom[2708] <= 8'b00000001;
font_rom[2709] <= 8'b00000000;
font_rom[2710] <= 8'b00000001;
font_rom[2711] <= 8'b00000000;
font_rom[2712] <= 8'b00000001;
font_rom[2713] <= 8'b00000000;
font_rom[2714] <= 8'b00000000;
font_rom[2715] <= 8'b00000000;
font_rom[2716] <= 8'b00000000;
font_rom[2717] <= 8'b00000000;
font_rom[2718] <= 8'b00000000;
font_rom[2719] <= 8'b00000000;
//ASCII 0x55 'U'
font_rom[2720] <= 8'b00000000;
font_rom[2721] <= 8'b00000000;
font_rom[2722] <= 8'b00000000;
font_rom[2723] <= 8'b00000000;
font_rom[2724] <= 8'b00000000;
font_rom[2725] <= 8'b00000000;
font_rom[2726] <= 8'b00000000;
font_rom[2727] <= 8'b00000000;
font_rom[2728] <= 8'b00000000;
font_rom[2729] <= 8'b00000000;
font_rom[2730] <= 8'b00001100;
font_rom[2731] <= 8'b00100000;
font_rom[2732] <= 8'b00001100;
font_rom[2733] <= 8'b00100000;
font_rom[2734] <= 8'b00001100;
font_rom[2735] <= 8'b00100000;
font_rom[2736] <= 8'b00001100;
font_rom[2737] <= 8'b01100000;
font_rom[2738] <= 8'b00001100;
font_rom[2739] <= 8'b01100000;
font_rom[2740] <= 8'b00001100;
font_rom[2741] <= 8'b01100000;
font_rom[2742] <= 8'b00000100;
font_rom[2743] <= 8'b01100000;
font_rom[2744] <= 8'b00000111;
font_rom[2745] <= 8'b11000000;
font_rom[2746] <= 8'b00000000;
font_rom[2747] <= 8'b00000000;
font_rom[2748] <= 8'b00000000;
font_rom[2749] <= 8'b00000000;
font_rom[2750] <= 8'b00000000;
font_rom[2751] <= 8'b00000000;
//ASCII 0x56 'V'
font_rom[2752] <= 8'b00000000;
font_rom[2753] <= 8'b00000000;
font_rom[2754] <= 8'b00000000;
font_rom[2755] <= 8'b00000000;
font_rom[2756] <= 8'b00000000;
font_rom[2757] <= 8'b00000000;
font_rom[2758] <= 8'b00000000;
font_rom[2759] <= 8'b00000000;
font_rom[2760] <= 8'b00000000;
font_rom[2761] <= 8'b00000000;
font_rom[2762] <= 8'b00001100;
font_rom[2763] <= 8'b01100000;
font_rom[2764] <= 8'b00001100;
font_rom[2765] <= 8'b01100000;
font_rom[2766] <= 8'b00000100;
font_rom[2767] <= 8'b11000000;
font_rom[2768] <= 8'b00000110;
font_rom[2769] <= 8'b11000000;
font_rom[2770] <= 8'b00000110;
font_rom[2771] <= 8'b11000000;
font_rom[2772] <= 8'b00000111;
font_rom[2773] <= 8'b10000000;
font_rom[2774] <= 8'b00000011;
font_rom[2775] <= 8'b10000000;
font_rom[2776] <= 8'b00000011;
font_rom[2777] <= 8'b00000000;
font_rom[2778] <= 8'b00000000;
font_rom[2779] <= 8'b00000000;
font_rom[2780] <= 8'b00000000;
font_rom[2781] <= 8'b00000000;
font_rom[2782] <= 8'b00000000;
font_rom[2783] <= 8'b00000000;
//ASCII 0x57 'W'
font_rom[2784] <= 8'b00000000;
font_rom[2785] <= 8'b00000000;
font_rom[2786] <= 8'b00000000;
font_rom[2787] <= 8'b00000000;
font_rom[2788] <= 8'b00000000;
font_rom[2789] <= 8'b00000000;
font_rom[2790] <= 8'b00000000;
font_rom[2791] <= 8'b00000000;
font_rom[2792] <= 8'b00000000;
font_rom[2793] <= 8'b00000000;
font_rom[2794] <= 8'b00110001;
font_rom[2795] <= 8'b10011000;
font_rom[2796] <= 8'b00110011;
font_rom[2797] <= 8'b10011000;
font_rom[2798] <= 8'b00011011;
font_rom[2799] <= 8'b10011000;
font_rom[2800] <= 8'b00011011;
font_rom[2801] <= 8'b10110000;
font_rom[2802] <= 8'b00011110;
font_rom[2803] <= 8'b10110000;
font_rom[2804] <= 8'b00011110;
font_rom[2805] <= 8'b11100000;
font_rom[2806] <= 8'b00001100;
font_rom[2807] <= 8'b11100000;
font_rom[2808] <= 8'b00001100;
font_rom[2809] <= 8'b11100000;
font_rom[2810] <= 8'b00000000;
font_rom[2811] <= 8'b00000000;
font_rom[2812] <= 8'b00000000;
font_rom[2813] <= 8'b00000000;
font_rom[2814] <= 8'b00000000;
font_rom[2815] <= 8'b00000000;
//ASCII 0x58 'X'
font_rom[2816] <= 8'b00000000;
font_rom[2817] <= 8'b00000000;
font_rom[2818] <= 8'b00000000;
font_rom[2819] <= 8'b00000000;
font_rom[2820] <= 8'b00000000;
font_rom[2821] <= 8'b00000000;
font_rom[2822] <= 8'b00000000;
font_rom[2823] <= 8'b00000000;
font_rom[2824] <= 8'b00000000;
font_rom[2825] <= 8'b00000000;
font_rom[2826] <= 8'b00001100;
font_rom[2827] <= 8'b00110000;
font_rom[2828] <= 8'b00000110;
font_rom[2829] <= 8'b01100000;
font_rom[2830] <= 8'b00000011;
font_rom[2831] <= 8'b11000000;
font_rom[2832] <= 8'b00000011;
font_rom[2833] <= 8'b10000000;
font_rom[2834] <= 8'b00000011;
font_rom[2835] <= 8'b10000000;
font_rom[2836] <= 8'b00000111;
font_rom[2837] <= 8'b11000000;
font_rom[2838] <= 8'b00001110;
font_rom[2839] <= 8'b01100000;
font_rom[2840] <= 8'b00001100;
font_rom[2841] <= 8'b01110000;
font_rom[2842] <= 8'b00000000;
font_rom[2843] <= 8'b00000000;
font_rom[2844] <= 8'b00000000;
font_rom[2845] <= 8'b00000000;
font_rom[2846] <= 8'b00000000;
font_rom[2847] <= 8'b00000000;
//ASCII 0x59 'Y'
font_rom[2848] <= 8'b00000000;
font_rom[2849] <= 8'b00000000;
font_rom[2850] <= 8'b00000000;
font_rom[2851] <= 8'b00000000;
font_rom[2852] <= 8'b00000000;
font_rom[2853] <= 8'b00000000;
font_rom[2854] <= 8'b00000000;
font_rom[2855] <= 8'b00000000;
font_rom[2856] <= 8'b00000000;
font_rom[2857] <= 8'b00000000;
font_rom[2858] <= 8'b00011000;
font_rom[2859] <= 8'b01100000;
font_rom[2860] <= 8'b00001100;
font_rom[2861] <= 8'b11000000;
font_rom[2862] <= 8'b00000110;
font_rom[2863] <= 8'b11000000;
font_rom[2864] <= 8'b00000111;
font_rom[2865] <= 8'b10000000;
font_rom[2866] <= 8'b00000011;
font_rom[2867] <= 8'b10000000;
font_rom[2868] <= 8'b00000011;
font_rom[2869] <= 8'b10000000;
font_rom[2870] <= 8'b00000011;
font_rom[2871] <= 8'b00000000;
font_rom[2872] <= 8'b00000110;
font_rom[2873] <= 8'b00000000;
font_rom[2874] <= 8'b00000000;
font_rom[2875] <= 8'b00000000;
font_rom[2876] <= 8'b00000000;
font_rom[2877] <= 8'b00000000;
font_rom[2878] <= 8'b00000000;
font_rom[2879] <= 8'b00000000;
//ASCII 0x5A 'Z'
font_rom[2880] <= 8'b00000000;
font_rom[2881] <= 8'b00000000;
font_rom[2882] <= 8'b00000000;
font_rom[2883] <= 8'b00000000;
font_rom[2884] <= 8'b00000000;
font_rom[2885] <= 8'b00000000;
font_rom[2886] <= 8'b00000000;
font_rom[2887] <= 8'b00000000;
font_rom[2888] <= 8'b00000000;
font_rom[2889] <= 8'b00000000;
font_rom[2890] <= 8'b00001111;
font_rom[2891] <= 8'b11110000;
font_rom[2892] <= 8'b00000000;
font_rom[2893] <= 8'b11100000;
font_rom[2894] <= 8'b00000001;
font_rom[2895] <= 8'b10000000;
font_rom[2896] <= 8'b00000011;
font_rom[2897] <= 8'b00000000;
font_rom[2898] <= 8'b00000011;
font_rom[2899] <= 8'b00000000;
font_rom[2900] <= 8'b00000110;
font_rom[2901] <= 8'b00000000;
font_rom[2902] <= 8'b00001100;
font_rom[2903] <= 8'b00000000;
font_rom[2904] <= 8'b00001111;
font_rom[2905] <= 8'b11110000;
font_rom[2906] <= 8'b00000000;
font_rom[2907] <= 8'b00000000;
font_rom[2908] <= 8'b00000000;
font_rom[2909] <= 8'b00000000;
font_rom[2910] <= 8'b00000000;
font_rom[2911] <= 8'b00000000;
//ASCII 0x5B '['
font_rom[2912] <= 8'b00000000;
font_rom[2913] <= 8'b00000000;
font_rom[2914] <= 8'b00000000;
font_rom[2915] <= 8'b00000000;
font_rom[2916] <= 8'b00000000;
font_rom[2917] <= 8'b00000000;
font_rom[2918] <= 8'b00000000;
font_rom[2919] <= 8'b00000000;
font_rom[2920] <= 8'b00000011;
font_rom[2921] <= 8'b11000000;
font_rom[2922] <= 8'b00000011;
font_rom[2923] <= 8'b00000000;
font_rom[2924] <= 8'b00000011;
font_rom[2925] <= 8'b00000000;
font_rom[2926] <= 8'b00000011;
font_rom[2927] <= 8'b00000000;
font_rom[2928] <= 8'b00000011;
font_rom[2929] <= 8'b00000000;
font_rom[2930] <= 8'b00000011;
font_rom[2931] <= 8'b00000000;
font_rom[2932] <= 8'b00000011;
font_rom[2933] <= 8'b00000000;
font_rom[2934] <= 8'b00000011;
font_rom[2935] <= 8'b00000000;
font_rom[2936] <= 8'b00000011;
font_rom[2937] <= 8'b00000000;
font_rom[2938] <= 8'b00000011;
font_rom[2939] <= 8'b00000000;
font_rom[2940] <= 8'b00000011;
font_rom[2941] <= 8'b11000000;
font_rom[2942] <= 8'b00000000;
font_rom[2943] <= 8'b00000000;
//ASCII 0x5C '\'
font_rom[2944] <= 8'b00000000;
font_rom[2945] <= 8'b00000000;
font_rom[2946] <= 8'b00000000;
font_rom[2947] <= 8'b00000000;
font_rom[2948] <= 8'b00000000;
font_rom[2949] <= 8'b00000000;
font_rom[2950] <= 8'b00000000;
font_rom[2951] <= 8'b00000000;
font_rom[2952] <= 8'b00000000;
font_rom[2953] <= 8'b00000000;
font_rom[2954] <= 8'b00000011;
font_rom[2955] <= 8'b00000000;
font_rom[2956] <= 8'b00000001;
font_rom[2957] <= 8'b10000000;
font_rom[2958] <= 8'b00000001;
font_rom[2959] <= 8'b10000000;
font_rom[2960] <= 8'b00000000;
font_rom[2961] <= 8'b11000000;
font_rom[2962] <= 8'b00000000;
font_rom[2963] <= 8'b11000000;
font_rom[2964] <= 8'b00000000;
font_rom[2965] <= 8'b11000000;
font_rom[2966] <= 8'b00000000;
font_rom[2967] <= 8'b01100000;
font_rom[2968] <= 8'b00000000;
font_rom[2969] <= 8'b01100000;
font_rom[2970] <= 8'b00000000;
font_rom[2971] <= 8'b00110000;
font_rom[2972] <= 8'b00000000;
font_rom[2973] <= 8'b00000000;
font_rom[2974] <= 8'b00000000;
font_rom[2975] <= 8'b00000000;
//ASCII 0x5D ']'
font_rom[2976] <= 8'b00000000;
font_rom[2977] <= 8'b00000000;
font_rom[2978] <= 8'b00000000;
font_rom[2979] <= 8'b00000000;
font_rom[2980] <= 8'b00000000;
font_rom[2981] <= 8'b00000000;
font_rom[2982] <= 8'b00000000;
font_rom[2983] <= 8'b00000000;
font_rom[2984] <= 8'b00000011;
font_rom[2985] <= 8'b11000000;
font_rom[2986] <= 8'b00000000;
font_rom[2987] <= 8'b11000000;
font_rom[2988] <= 8'b00000000;
font_rom[2989] <= 8'b11000000;
font_rom[2990] <= 8'b00000000;
font_rom[2991] <= 8'b11000000;
font_rom[2992] <= 8'b00000000;
font_rom[2993] <= 8'b11000000;
font_rom[2994] <= 8'b00000000;
font_rom[2995] <= 8'b11000000;
font_rom[2996] <= 8'b00000000;
font_rom[2997] <= 8'b11000000;
font_rom[2998] <= 8'b00000000;
font_rom[2999] <= 8'b11000000;
font_rom[3000] <= 8'b00000000;
font_rom[3001] <= 8'b11000000;
font_rom[3002] <= 8'b00000000;
font_rom[3003] <= 8'b11000000;
font_rom[3004] <= 8'b00000011;
font_rom[3005] <= 8'b11000000;
font_rom[3006] <= 8'b00000000;
font_rom[3007] <= 8'b00000000;
//ASCII 0x5E '^'
font_rom[3008] <= 8'b00000000;
font_rom[3009] <= 8'b00000000;
font_rom[3010] <= 8'b00000000;
font_rom[3011] <= 8'b00000000;
font_rom[3012] <= 8'b00000000;
font_rom[3013] <= 8'b00000000;
font_rom[3014] <= 8'b00000000;
font_rom[3015] <= 8'b00000000;
font_rom[3016] <= 8'b00000000;
font_rom[3017] <= 8'b11000000;
font_rom[3018] <= 8'b00000001;
font_rom[3019] <= 8'b11100000;
font_rom[3020] <= 8'b00000011;
font_rom[3021] <= 8'b00110000;
font_rom[3022] <= 8'b00000000;
font_rom[3023] <= 8'b00000000;
font_rom[3024] <= 8'b00000000;
font_rom[3025] <= 8'b00000000;
font_rom[3026] <= 8'b00000000;
font_rom[3027] <= 8'b00000000;
font_rom[3028] <= 8'b00000000;
font_rom[3029] <= 8'b00000000;
font_rom[3030] <= 8'b00000000;
font_rom[3031] <= 8'b00000000;
font_rom[3032] <= 8'b00000000;
font_rom[3033] <= 8'b00000000;
font_rom[3034] <= 8'b00000000;
font_rom[3035] <= 8'b00000000;
font_rom[3036] <= 8'b00000000;
font_rom[3037] <= 8'b00000000;
font_rom[3038] <= 8'b00000000;
font_rom[3039] <= 8'b00000000;
//ASCII 0x5F '_'
font_rom[3040] <= 8'b00000000;
font_rom[3041] <= 8'b00000000;
font_rom[3042] <= 8'b00000000;
font_rom[3043] <= 8'b00000000;
font_rom[3044] <= 8'b00000000;
font_rom[3045] <= 8'b00000000;
font_rom[3046] <= 8'b00000000;
font_rom[3047] <= 8'b00000000;
font_rom[3048] <= 8'b00000000;
font_rom[3049] <= 8'b00000000;
font_rom[3050] <= 8'b00000000;
font_rom[3051] <= 8'b00000000;
font_rom[3052] <= 8'b00000000;
font_rom[3053] <= 8'b00000000;
font_rom[3054] <= 8'b00000000;
font_rom[3055] <= 8'b00000000;
font_rom[3056] <= 8'b00000000;
font_rom[3057] <= 8'b00000000;
font_rom[3058] <= 8'b00000000;
font_rom[3059] <= 8'b00000000;
font_rom[3060] <= 8'b00000000;
font_rom[3061] <= 8'b00000000;
font_rom[3062] <= 8'b00000000;
font_rom[3063] <= 8'b00000000;
font_rom[3064] <= 8'b00000000;
font_rom[3065] <= 8'b00000000;
font_rom[3066] <= 8'b00000000;
font_rom[3067] <= 8'b00000000;
font_rom[3068] <= 8'b00011111;
font_rom[3069] <= 8'b11100000;
font_rom[3070] <= 8'b00000000;
font_rom[3071] <= 8'b00000000;
//ASCII 0x60 '`'
font_rom[3072] <= 8'b00000000;
font_rom[3073] <= 8'b00000000;
font_rom[3074] <= 8'b00000000;
font_rom[3075] <= 8'b00000000;
font_rom[3076] <= 8'b00000000;
font_rom[3077] <= 8'b00000000;
font_rom[3078] <= 8'b00000000;
font_rom[3079] <= 8'b00000000;
font_rom[3080] <= 8'b00000110;
font_rom[3081] <= 8'b00000000;
font_rom[3082] <= 8'b00000011;
font_rom[3083] <= 8'b00000000;
font_rom[3084] <= 8'b00000000;
font_rom[3085] <= 8'b00000000;
font_rom[3086] <= 8'b00000000;
font_rom[3087] <= 8'b00000000;
font_rom[3088] <= 8'b00000000;
font_rom[3089] <= 8'b00000000;
font_rom[3090] <= 8'b00000000;
font_rom[3091] <= 8'b00000000;
font_rom[3092] <= 8'b00000000;
font_rom[3093] <= 8'b00000000;
font_rom[3094] <= 8'b00000000;
font_rom[3095] <= 8'b00000000;
font_rom[3096] <= 8'b00000000;
font_rom[3097] <= 8'b00000000;
font_rom[3098] <= 8'b00000000;
font_rom[3099] <= 8'b00000000;
font_rom[3100] <= 8'b00000000;
font_rom[3101] <= 8'b00000000;
font_rom[3102] <= 8'b00000000;
font_rom[3103] <= 8'b00000000;
//ASCII 0x61 'a'
font_rom[3104] <= 8'b00000000;
font_rom[3105] <= 8'b00000000;
font_rom[3106] <= 8'b00000000;
font_rom[3107] <= 8'b00000000;
font_rom[3108] <= 8'b00000000;
font_rom[3109] <= 8'b00000000;
font_rom[3110] <= 8'b00000000;
font_rom[3111] <= 8'b00000000;
font_rom[3112] <= 8'b00000000;
font_rom[3113] <= 8'b00000000;
font_rom[3114] <= 8'b00000000;
font_rom[3115] <= 8'b00000000;
font_rom[3116] <= 8'b00000000;
font_rom[3117] <= 8'b00000000;
font_rom[3118] <= 8'b00000011;
font_rom[3119] <= 8'b11000000;
font_rom[3120] <= 8'b00000110;
font_rom[3121] <= 8'b11000000;
font_rom[3122] <= 8'b00000110;
font_rom[3123] <= 8'b11000000;
font_rom[3124] <= 8'b00000100;
font_rom[3125] <= 8'b11000000;
font_rom[3126] <= 8'b00000110;
font_rom[3127] <= 8'b11000000;
font_rom[3128] <= 8'b00000111;
font_rom[3129] <= 8'b11100000;
font_rom[3130] <= 8'b00000000;
font_rom[3131] <= 8'b00000000;
font_rom[3132] <= 8'b00000000;
font_rom[3133] <= 8'b00000000;
font_rom[3134] <= 8'b00000000;
font_rom[3135] <= 8'b00000000;
//ASCII 0x62 'b'
font_rom[3136] <= 8'b00000000;
font_rom[3137] <= 8'b00000000;
font_rom[3138] <= 8'b00000000;
font_rom[3139] <= 8'b00000000;
font_rom[3140] <= 8'b00000000;
font_rom[3141] <= 8'b00000000;
font_rom[3142] <= 8'b00000000;
font_rom[3143] <= 8'b00000000;
font_rom[3144] <= 8'b00000110;
font_rom[3145] <= 8'b00000000;
font_rom[3146] <= 8'b00000110;
font_rom[3147] <= 8'b00000000;
font_rom[3148] <= 8'b00000110;
font_rom[3149] <= 8'b00000000;
font_rom[3150] <= 8'b00000111;
font_rom[3151] <= 8'b11000000;
font_rom[3152] <= 8'b00000110;
font_rom[3153] <= 8'b01000000;
font_rom[3154] <= 8'b00000110;
font_rom[3155] <= 8'b01100000;
font_rom[3156] <= 8'b00000110;
font_rom[3157] <= 8'b01100000;
font_rom[3158] <= 8'b00000110;
font_rom[3159] <= 8'b11000000;
font_rom[3160] <= 8'b00000111;
font_rom[3161] <= 8'b11000000;
font_rom[3162] <= 8'b00000000;
font_rom[3163] <= 8'b00000000;
font_rom[3164] <= 8'b00000000;
font_rom[3165] <= 8'b00000000;
font_rom[3166] <= 8'b00000000;
font_rom[3167] <= 8'b00000000;
//ASCII 0x63 'c'
font_rom[3168] <= 8'b00000000;
font_rom[3169] <= 8'b00000000;
font_rom[3170] <= 8'b00000000;
font_rom[3171] <= 8'b00000000;
font_rom[3172] <= 8'b00000000;
font_rom[3173] <= 8'b00000000;
font_rom[3174] <= 8'b00000000;
font_rom[3175] <= 8'b00000000;
font_rom[3176] <= 8'b00000000;
font_rom[3177] <= 8'b00000000;
font_rom[3178] <= 8'b00000000;
font_rom[3179] <= 8'b00000000;
font_rom[3180] <= 8'b00000000;
font_rom[3181] <= 8'b00000000;
font_rom[3182] <= 8'b00000001;
font_rom[3183] <= 8'b11000000;
font_rom[3184] <= 8'b00000011;
font_rom[3185] <= 8'b01100000;
font_rom[3186] <= 8'b00000110;
font_rom[3187] <= 8'b00000000;
font_rom[3188] <= 8'b00000110;
font_rom[3189] <= 8'b00000000;
font_rom[3190] <= 8'b00000110;
font_rom[3191] <= 8'b01100000;
font_rom[3192] <= 8'b00000011;
font_rom[3193] <= 8'b11000000;
font_rom[3194] <= 8'b00000000;
font_rom[3195] <= 8'b00000000;
font_rom[3196] <= 8'b00000000;
font_rom[3197] <= 8'b00000000;
font_rom[3198] <= 8'b00000000;
font_rom[3199] <= 8'b00000000;
//ASCII 0x64 'd'
font_rom[3200] <= 8'b00000000;
font_rom[3201] <= 8'b00000000;
font_rom[3202] <= 8'b00000000;
font_rom[3203] <= 8'b00000000;
font_rom[3204] <= 8'b00000000;
font_rom[3205] <= 8'b00000000;
font_rom[3206] <= 8'b00000000;
font_rom[3207] <= 8'b00000000;
font_rom[3208] <= 8'b00000000;
font_rom[3209] <= 8'b01100000;
font_rom[3210] <= 8'b00000000;
font_rom[3211] <= 8'b01100000;
font_rom[3212] <= 8'b00000000;
font_rom[3213] <= 8'b01000000;
font_rom[3214] <= 8'b00000011;
font_rom[3215] <= 8'b11000000;
font_rom[3216] <= 8'b00000110;
font_rom[3217] <= 8'b11000000;
font_rom[3218] <= 8'b00000110;
font_rom[3219] <= 8'b01000000;
font_rom[3220] <= 8'b00000110;
font_rom[3221] <= 8'b01000000;
font_rom[3222] <= 8'b00000110;
font_rom[3223] <= 8'b11000000;
font_rom[3224] <= 8'b00000011;
font_rom[3225] <= 8'b11100000;
font_rom[3226] <= 8'b00000000;
font_rom[3227] <= 8'b00000000;
font_rom[3228] <= 8'b00000000;
font_rom[3229] <= 8'b00000000;
font_rom[3230] <= 8'b00000000;
font_rom[3231] <= 8'b00000000;
//ASCII 0x65 'e'
font_rom[3232] <= 8'b00000000;
font_rom[3233] <= 8'b00000000;
font_rom[3234] <= 8'b00000000;
font_rom[3235] <= 8'b00000000;
font_rom[3236] <= 8'b00000000;
font_rom[3237] <= 8'b00000000;
font_rom[3238] <= 8'b00000000;
font_rom[3239] <= 8'b00000000;
font_rom[3240] <= 8'b00000000;
font_rom[3241] <= 8'b00000000;
font_rom[3242] <= 8'b00000000;
font_rom[3243] <= 8'b00000000;
font_rom[3244] <= 8'b00000000;
font_rom[3245] <= 8'b00000000;
font_rom[3246] <= 8'b00000011;
font_rom[3247] <= 8'b11000000;
font_rom[3248] <= 8'b00000110;
font_rom[3249] <= 8'b01000000;
font_rom[3250] <= 8'b00000111;
font_rom[3251] <= 8'b11000000;
font_rom[3252] <= 8'b00000111;
font_rom[3253] <= 8'b00000000;
font_rom[3254] <= 8'b00000110;
font_rom[3255] <= 8'b01100000;
font_rom[3256] <= 8'b00000011;
font_rom[3257] <= 8'b11000000;
font_rom[3258] <= 8'b00000000;
font_rom[3259] <= 8'b00000000;
font_rom[3260] <= 8'b00000000;
font_rom[3261] <= 8'b00000000;
font_rom[3262] <= 8'b00000000;
font_rom[3263] <= 8'b00000000;
//ASCII 0x66 'f'
font_rom[3264] <= 8'b00000000;
font_rom[3265] <= 8'b00000000;
font_rom[3266] <= 8'b00000000;
font_rom[3267] <= 8'b00000000;
font_rom[3268] <= 8'b00000000;
font_rom[3269] <= 8'b00000000;
font_rom[3270] <= 8'b00000000;
font_rom[3271] <= 8'b00000000;
font_rom[3272] <= 8'b00000001;
font_rom[3273] <= 8'b11000000;
font_rom[3274] <= 8'b00000001;
font_rom[3275] <= 8'b00000000;
font_rom[3276] <= 8'b00000011;
font_rom[3277] <= 8'b00000000;
font_rom[3278] <= 8'b00000111;
font_rom[3279] <= 8'b11000000;
font_rom[3280] <= 8'b00000011;
font_rom[3281] <= 8'b00000000;
font_rom[3282] <= 8'b00000011;
font_rom[3283] <= 8'b00000000;
font_rom[3284] <= 8'b00000011;
font_rom[3285] <= 8'b00000000;
font_rom[3286] <= 8'b00000011;
font_rom[3287] <= 8'b00000000;
font_rom[3288] <= 8'b00000011;
font_rom[3289] <= 8'b00000000;
font_rom[3290] <= 8'b00000000;
font_rom[3291] <= 8'b00000000;
font_rom[3292] <= 8'b00000000;
font_rom[3293] <= 8'b00000000;
font_rom[3294] <= 8'b00000000;
font_rom[3295] <= 8'b00000000;
//ASCII 0x67 'g'
font_rom[3296] <= 8'b00000000;
font_rom[3297] <= 8'b00000000;
font_rom[3298] <= 8'b00000000;
font_rom[3299] <= 8'b00000000;
font_rom[3300] <= 8'b00000000;
font_rom[3301] <= 8'b00000000;
font_rom[3302] <= 8'b00000000;
font_rom[3303] <= 8'b00000000;
font_rom[3304] <= 8'b00000000;
font_rom[3305] <= 8'b00000000;
font_rom[3306] <= 8'b00000000;
font_rom[3307] <= 8'b00000000;
font_rom[3308] <= 8'b00000000;
font_rom[3309] <= 8'b00000000;
font_rom[3310] <= 8'b00000011;
font_rom[3311] <= 8'b11000000;
font_rom[3312] <= 8'b00000110;
font_rom[3313] <= 8'b01100000;
font_rom[3314] <= 8'b00000110;
font_rom[3315] <= 8'b01100000;
font_rom[3316] <= 8'b00000100;
font_rom[3317] <= 8'b11000000;
font_rom[3318] <= 8'b00000110;
font_rom[3319] <= 8'b11000000;
font_rom[3320] <= 8'b00000111;
font_rom[3321] <= 8'b11000000;
font_rom[3322] <= 8'b00000000;
font_rom[3323] <= 8'b11000000;
font_rom[3324] <= 8'b00000000;
font_rom[3325] <= 8'b11000000;
font_rom[3326] <= 8'b00000111;
font_rom[3327] <= 8'b10000000;
//ASCII 0x68 'h'
font_rom[3328] <= 8'b00000000;
font_rom[3329] <= 8'b00000000;
font_rom[3330] <= 8'b00000000;
font_rom[3331] <= 8'b00000000;
font_rom[3332] <= 8'b00000000;
font_rom[3333] <= 8'b00000000;
font_rom[3334] <= 8'b00000000;
font_rom[3335] <= 8'b00000000;
font_rom[3336] <= 8'b00000110;
font_rom[3337] <= 8'b00000000;
font_rom[3338] <= 8'b00000110;
font_rom[3339] <= 8'b00000000;
font_rom[3340] <= 8'b00000110;
font_rom[3341] <= 8'b00000000;
font_rom[3342] <= 8'b00000111;
font_rom[3343] <= 8'b11000000;
font_rom[3344] <= 8'b00000111;
font_rom[3345] <= 8'b11000000;
font_rom[3346] <= 8'b00000110;
font_rom[3347] <= 8'b11000000;
font_rom[3348] <= 8'b00000110;
font_rom[3349] <= 8'b11000000;
font_rom[3350] <= 8'b00000110;
font_rom[3351] <= 8'b11000000;
font_rom[3352] <= 8'b00000110;
font_rom[3353] <= 8'b01100000;
font_rom[3354] <= 8'b00000000;
font_rom[3355] <= 8'b00000000;
font_rom[3356] <= 8'b00000000;
font_rom[3357] <= 8'b00000000;
font_rom[3358] <= 8'b00000000;
font_rom[3359] <= 8'b00000000;
//ASCII 0x69 'i'
font_rom[3360] <= 8'b00000000;
font_rom[3361] <= 8'b00000000;
font_rom[3362] <= 8'b00000000;
font_rom[3363] <= 8'b00000000;
font_rom[3364] <= 8'b00000000;
font_rom[3365] <= 8'b00000000;
font_rom[3366] <= 8'b00000000;
font_rom[3367] <= 8'b00000000;
font_rom[3368] <= 8'b00000000;
font_rom[3369] <= 8'b00000000;
font_rom[3370] <= 8'b00000001;
font_rom[3371] <= 8'b10000000;
font_rom[3372] <= 8'b00000000;
font_rom[3373] <= 8'b00000000;
font_rom[3374] <= 8'b00000001;
font_rom[3375] <= 8'b10000000;
font_rom[3376] <= 8'b00000001;
font_rom[3377] <= 8'b10000000;
font_rom[3378] <= 8'b00000001;
font_rom[3379] <= 8'b10000000;
font_rom[3380] <= 8'b00000001;
font_rom[3381] <= 8'b10000000;
font_rom[3382] <= 8'b00000001;
font_rom[3383] <= 8'b10000000;
font_rom[3384] <= 8'b00000001;
font_rom[3385] <= 8'b10000000;
font_rom[3386] <= 8'b00000000;
font_rom[3387] <= 8'b00000000;
font_rom[3388] <= 8'b00000000;
font_rom[3389] <= 8'b00000000;
font_rom[3390] <= 8'b00000000;
font_rom[3391] <= 8'b00000000;
//ASCII 0x6A 'j'
font_rom[3392] <= 8'b00000000;
font_rom[3393] <= 8'b00000000;
font_rom[3394] <= 8'b00000000;
font_rom[3395] <= 8'b00000000;
font_rom[3396] <= 8'b00000000;
font_rom[3397] <= 8'b00000000;
font_rom[3398] <= 8'b00000000;
font_rom[3399] <= 8'b00000000;
font_rom[3400] <= 8'b00000000;
font_rom[3401] <= 8'b00000000;
font_rom[3402] <= 8'b00000001;
font_rom[3403] <= 8'b10000000;
font_rom[3404] <= 8'b00000000;
font_rom[3405] <= 8'b00000000;
font_rom[3406] <= 8'b00000001;
font_rom[3407] <= 8'b10000000;
font_rom[3408] <= 8'b00000001;
font_rom[3409] <= 8'b10000000;
font_rom[3410] <= 8'b00000001;
font_rom[3411] <= 8'b10000000;
font_rom[3412] <= 8'b00000001;
font_rom[3413] <= 8'b10000000;
font_rom[3414] <= 8'b00000001;
font_rom[3415] <= 8'b10000000;
font_rom[3416] <= 8'b00000001;
font_rom[3417] <= 8'b10000000;
font_rom[3418] <= 8'b00000001;
font_rom[3419] <= 8'b10000000;
font_rom[3420] <= 8'b00000111;
font_rom[3421] <= 8'b10000000;
font_rom[3422] <= 8'b00000011;
font_rom[3423] <= 8'b10000000;
//ASCII 0x6B 'k'
font_rom[3424] <= 8'b00000000;
font_rom[3425] <= 8'b00000000;
font_rom[3426] <= 8'b00000000;
font_rom[3427] <= 8'b00000000;
font_rom[3428] <= 8'b00000000;
font_rom[3429] <= 8'b00000000;
font_rom[3430] <= 8'b00000000;
font_rom[3431] <= 8'b00000000;
font_rom[3432] <= 8'b00000110;
font_rom[3433] <= 8'b00000000;
font_rom[3434] <= 8'b00000110;
font_rom[3435] <= 8'b00000000;
font_rom[3436] <= 8'b00000110;
font_rom[3437] <= 8'b00000000;
font_rom[3438] <= 8'b00000110;
font_rom[3439] <= 8'b11100000;
font_rom[3440] <= 8'b00000110;
font_rom[3441] <= 8'b11000000;
font_rom[3442] <= 8'b00000111;
font_rom[3443] <= 8'b10000000;
font_rom[3444] <= 8'b00000111;
font_rom[3445] <= 8'b11000000;
font_rom[3446] <= 8'b00000110;
font_rom[3447] <= 8'b11000000;
font_rom[3448] <= 8'b00000110;
font_rom[3449] <= 8'b01100000;
font_rom[3450] <= 8'b00000000;
font_rom[3451] <= 8'b00000000;
font_rom[3452] <= 8'b00000000;
font_rom[3453] <= 8'b00000000;
font_rom[3454] <= 8'b00000000;
font_rom[3455] <= 8'b00000000;
//ASCII 0x6C 'l'
font_rom[3456] <= 8'b00000000;
font_rom[3457] <= 8'b00000000;
font_rom[3458] <= 8'b00000000;
font_rom[3459] <= 8'b00000000;
font_rom[3460] <= 8'b00000000;
font_rom[3461] <= 8'b00000000;
font_rom[3462] <= 8'b00000000;
font_rom[3463] <= 8'b00000000;
font_rom[3464] <= 8'b00000011;
font_rom[3465] <= 8'b00000000;
font_rom[3466] <= 8'b00000011;
font_rom[3467] <= 8'b00000000;
font_rom[3468] <= 8'b00000011;
font_rom[3469] <= 8'b00000000;
font_rom[3470] <= 8'b00000011;
font_rom[3471] <= 8'b00000000;
font_rom[3472] <= 8'b00000011;
font_rom[3473] <= 8'b00000000;
font_rom[3474] <= 8'b00000011;
font_rom[3475] <= 8'b00000000;
font_rom[3476] <= 8'b00000011;
font_rom[3477] <= 8'b00000000;
font_rom[3478] <= 8'b00000011;
font_rom[3479] <= 8'b00000000;
font_rom[3480] <= 8'b00000011;
font_rom[3481] <= 8'b00000000;
font_rom[3482] <= 8'b00000000;
font_rom[3483] <= 8'b00000000;
font_rom[3484] <= 8'b00000000;
font_rom[3485] <= 8'b00000000;
font_rom[3486] <= 8'b00000000;
font_rom[3487] <= 8'b00000000;
//ASCII 0x6D 'm'
font_rom[3488] <= 8'b00000000;
font_rom[3489] <= 8'b00000000;
font_rom[3490] <= 8'b00000000;
font_rom[3491] <= 8'b00000000;
font_rom[3492] <= 8'b00000000;
font_rom[3493] <= 8'b00000000;
font_rom[3494] <= 8'b00000000;
font_rom[3495] <= 8'b00000000;
font_rom[3496] <= 8'b00000000;
font_rom[3497] <= 8'b00000000;
font_rom[3498] <= 8'b00000000;
font_rom[3499] <= 8'b00000000;
font_rom[3500] <= 8'b00000000;
font_rom[3501] <= 8'b00000000;
font_rom[3502] <= 8'b00001111;
font_rom[3503] <= 8'b11100000;
font_rom[3504] <= 8'b00001111;
font_rom[3505] <= 8'b11100000;
font_rom[3506] <= 8'b00001101;
font_rom[3507] <= 8'b11100000;
font_rom[3508] <= 8'b00001101;
font_rom[3509] <= 8'b10100000;
font_rom[3510] <= 8'b00001101;
font_rom[3511] <= 8'b10110000;
font_rom[3512] <= 8'b00001101;
font_rom[3513] <= 8'b10110000;
font_rom[3514] <= 8'b00000000;
font_rom[3515] <= 8'b00000000;
font_rom[3516] <= 8'b00000000;
font_rom[3517] <= 8'b00000000;
font_rom[3518] <= 8'b00000000;
font_rom[3519] <= 8'b00000000;
//ASCII 0x6E 'n'
font_rom[3520] <= 8'b00000000;
font_rom[3521] <= 8'b00000000;
font_rom[3522] <= 8'b00000000;
font_rom[3523] <= 8'b00000000;
font_rom[3524] <= 8'b00000000;
font_rom[3525] <= 8'b00000000;
font_rom[3526] <= 8'b00000000;
font_rom[3527] <= 8'b00000000;
font_rom[3528] <= 8'b00000000;
font_rom[3529] <= 8'b00000000;
font_rom[3530] <= 8'b00000000;
font_rom[3531] <= 8'b00000000;
font_rom[3532] <= 8'b00000000;
font_rom[3533] <= 8'b00000000;
font_rom[3534] <= 8'b00000111;
font_rom[3535] <= 8'b11000000;
font_rom[3536] <= 8'b00000111;
font_rom[3537] <= 8'b11000000;
font_rom[3538] <= 8'b00000110;
font_rom[3539] <= 8'b01100000;
font_rom[3540] <= 8'b00000110;
font_rom[3541] <= 8'b01100000;
font_rom[3542] <= 8'b00000110;
font_rom[3543] <= 8'b01100000;
font_rom[3544] <= 8'b00000110;
font_rom[3545] <= 8'b01100000;
font_rom[3546] <= 8'b00000000;
font_rom[3547] <= 8'b00000000;
font_rom[3548] <= 8'b00000000;
font_rom[3549] <= 8'b00000000;
font_rom[3550] <= 8'b00000000;
font_rom[3551] <= 8'b00000000;
//ASCII 0x6F 'o'
font_rom[3552] <= 8'b00000000;
font_rom[3553] <= 8'b00000000;
font_rom[3554] <= 8'b00000000;
font_rom[3555] <= 8'b00000000;
font_rom[3556] <= 8'b00000000;
font_rom[3557] <= 8'b00000000;
font_rom[3558] <= 8'b00000000;
font_rom[3559] <= 8'b00000000;
font_rom[3560] <= 8'b00000000;
font_rom[3561] <= 8'b00000000;
font_rom[3562] <= 8'b00000000;
font_rom[3563] <= 8'b00000000;
font_rom[3564] <= 8'b00000000;
font_rom[3565] <= 8'b00000000;
font_rom[3566] <= 8'b00000011;
font_rom[3567] <= 8'b11000000;
font_rom[3568] <= 8'b00000110;
font_rom[3569] <= 8'b11000000;
font_rom[3570] <= 8'b00000110;
font_rom[3571] <= 8'b01000000;
font_rom[3572] <= 8'b00000110;
font_rom[3573] <= 8'b01000000;
font_rom[3574] <= 8'b00000110;
font_rom[3575] <= 8'b11000000;
font_rom[3576] <= 8'b00000011;
font_rom[3577] <= 8'b10000000;
font_rom[3578] <= 8'b00000000;
font_rom[3579] <= 8'b00000000;
font_rom[3580] <= 8'b00000000;
font_rom[3581] <= 8'b00000000;
font_rom[3582] <= 8'b00000000;
font_rom[3583] <= 8'b00000000;
//ASCII 0x70 'p'
font_rom[3584] <= 8'b00000000;
font_rom[3585] <= 8'b00000000;
font_rom[3586] <= 8'b00000000;
font_rom[3587] <= 8'b00000000;
font_rom[3588] <= 8'b00000000;
font_rom[3589] <= 8'b00000000;
font_rom[3590] <= 8'b00000000;
font_rom[3591] <= 8'b00000000;
font_rom[3592] <= 8'b00000000;
font_rom[3593] <= 8'b00000000;
font_rom[3594] <= 8'b00000000;
font_rom[3595] <= 8'b00000000;
font_rom[3596] <= 8'b00000000;
font_rom[3597] <= 8'b00000000;
font_rom[3598] <= 8'b00000111;
font_rom[3599] <= 8'b11000000;
font_rom[3600] <= 8'b00000110;
font_rom[3601] <= 8'b11000000;
font_rom[3602] <= 8'b00000110;
font_rom[3603] <= 8'b01100000;
font_rom[3604] <= 8'b00000110;
font_rom[3605] <= 8'b01100000;
font_rom[3606] <= 8'b00000110;
font_rom[3607] <= 8'b11000000;
font_rom[3608] <= 8'b00000111;
font_rom[3609] <= 8'b11000000;
font_rom[3610] <= 8'b00000110;
font_rom[3611] <= 8'b00000000;
font_rom[3612] <= 8'b00000110;
font_rom[3613] <= 8'b00000000;
font_rom[3614] <= 8'b00000110;
font_rom[3615] <= 8'b00000000;
//ASCII 0x71 'q'
font_rom[3616] <= 8'b00000000;
font_rom[3617] <= 8'b00000000;
font_rom[3618] <= 8'b00000000;
font_rom[3619] <= 8'b00000000;
font_rom[3620] <= 8'b00000000;
font_rom[3621] <= 8'b00000000;
font_rom[3622] <= 8'b00000000;
font_rom[3623] <= 8'b00000000;
font_rom[3624] <= 8'b00000000;
font_rom[3625] <= 8'b00000000;
font_rom[3626] <= 8'b00000000;
font_rom[3627] <= 8'b00000000;
font_rom[3628] <= 8'b00000000;
font_rom[3629] <= 8'b00000000;
font_rom[3630] <= 8'b00000011;
font_rom[3631] <= 8'b11000000;
font_rom[3632] <= 8'b00000110;
font_rom[3633] <= 8'b11000000;
font_rom[3634] <= 8'b00000110;
font_rom[3635] <= 8'b11000000;
font_rom[3636] <= 8'b00000110;
font_rom[3637] <= 8'b11000000;
font_rom[3638] <= 8'b00000110;
font_rom[3639] <= 8'b11000000;
font_rom[3640] <= 8'b00000011;
font_rom[3641] <= 8'b11000000;
font_rom[3642] <= 8'b00000000;
font_rom[3643] <= 8'b11000000;
font_rom[3644] <= 8'b00000000;
font_rom[3645] <= 8'b11000000;
font_rom[3646] <= 8'b00000000;
font_rom[3647] <= 8'b11000000;
//ASCII 0x72 'r'
font_rom[3648] <= 8'b00000000;
font_rom[3649] <= 8'b00000000;
font_rom[3650] <= 8'b00000000;
font_rom[3651] <= 8'b00000000;
font_rom[3652] <= 8'b00000000;
font_rom[3653] <= 8'b00000000;
font_rom[3654] <= 8'b00000000;
font_rom[3655] <= 8'b00000000;
font_rom[3656] <= 8'b00000000;
font_rom[3657] <= 8'b00000000;
font_rom[3658] <= 8'b00000000;
font_rom[3659] <= 8'b00000000;
font_rom[3660] <= 8'b00000000;
font_rom[3661] <= 8'b00000000;
font_rom[3662] <= 8'b00000011;
font_rom[3663] <= 8'b11100000;
font_rom[3664] <= 8'b00000011;
font_rom[3665] <= 8'b01100000;
font_rom[3666] <= 8'b00000011;
font_rom[3667] <= 8'b00000000;
font_rom[3668] <= 8'b00000011;
font_rom[3669] <= 8'b00000000;
font_rom[3670] <= 8'b00000011;
font_rom[3671] <= 8'b00000000;
font_rom[3672] <= 8'b00000011;
font_rom[3673] <= 8'b00000000;
font_rom[3674] <= 8'b00000000;
font_rom[3675] <= 8'b00000000;
font_rom[3676] <= 8'b00000000;
font_rom[3677] <= 8'b00000000;
font_rom[3678] <= 8'b00000000;
font_rom[3679] <= 8'b00000000;
//ASCII 0x73 's'
font_rom[3680] <= 8'b00000000;
font_rom[3681] <= 8'b00000000;
font_rom[3682] <= 8'b00000000;
font_rom[3683] <= 8'b00000000;
font_rom[3684] <= 8'b00000000;
font_rom[3685] <= 8'b00000000;
font_rom[3686] <= 8'b00000000;
font_rom[3687] <= 8'b00000000;
font_rom[3688] <= 8'b00000000;
font_rom[3689] <= 8'b00000000;
font_rom[3690] <= 8'b00000000;
font_rom[3691] <= 8'b00000000;
font_rom[3692] <= 8'b00000000;
font_rom[3693] <= 8'b00000000;
font_rom[3694] <= 8'b00000000;
font_rom[3695] <= 8'b11100000;
font_rom[3696] <= 8'b00000011;
font_rom[3697] <= 8'b00000000;
font_rom[3698] <= 8'b00000011;
font_rom[3699] <= 8'b10000000;
font_rom[3700] <= 8'b00000000;
font_rom[3701] <= 8'b11000000;
font_rom[3702] <= 8'b00000000;
font_rom[3703] <= 8'b01100000;
font_rom[3704] <= 8'b00000111;
font_rom[3705] <= 8'b11000000;
font_rom[3706] <= 8'b00000000;
font_rom[3707] <= 8'b00000000;
font_rom[3708] <= 8'b00000000;
font_rom[3709] <= 8'b00000000;
font_rom[3710] <= 8'b00000000;
font_rom[3711] <= 8'b00000000;
//ASCII 0x74 't'
font_rom[3712] <= 8'b00000000;
font_rom[3713] <= 8'b00000000;
font_rom[3714] <= 8'b00000000;
font_rom[3715] <= 8'b00000000;
font_rom[3716] <= 8'b00000000;
font_rom[3717] <= 8'b00000000;
font_rom[3718] <= 8'b00000000;
font_rom[3719] <= 8'b00000000;
font_rom[3720] <= 8'b00000000;
font_rom[3721] <= 8'b00000000;
font_rom[3722] <= 8'b00000001;
font_rom[3723] <= 8'b10000000;
font_rom[3724] <= 8'b00000001;
font_rom[3725] <= 8'b10000000;
font_rom[3726] <= 8'b00000111;
font_rom[3727] <= 8'b11000000;
font_rom[3728] <= 8'b00000001;
font_rom[3729] <= 8'b10000000;
font_rom[3730] <= 8'b00000001;
font_rom[3731] <= 8'b10000000;
font_rom[3732] <= 8'b00000001;
font_rom[3733] <= 8'b10000000;
font_rom[3734] <= 8'b00000001;
font_rom[3735] <= 8'b10000000;
font_rom[3736] <= 8'b00000001;
font_rom[3737] <= 8'b10000000;
font_rom[3738] <= 8'b00000000;
font_rom[3739] <= 8'b00000000;
font_rom[3740] <= 8'b00000000;
font_rom[3741] <= 8'b00000000;
font_rom[3742] <= 8'b00000000;
font_rom[3743] <= 8'b00000000;
//ASCII 0x75 'u'
font_rom[3744] <= 8'b00000000;
font_rom[3745] <= 8'b00000000;
font_rom[3746] <= 8'b00000000;
font_rom[3747] <= 8'b00000000;
font_rom[3748] <= 8'b00000000;
font_rom[3749] <= 8'b00000000;
font_rom[3750] <= 8'b00000000;
font_rom[3751] <= 8'b00000000;
font_rom[3752] <= 8'b00000000;
font_rom[3753] <= 8'b00000000;
font_rom[3754] <= 8'b00000000;
font_rom[3755] <= 8'b00000000;
font_rom[3756] <= 8'b00000000;
font_rom[3757] <= 8'b00000000;
font_rom[3758] <= 8'b00000110;
font_rom[3759] <= 8'b01000000;
font_rom[3760] <= 8'b00000110;
font_rom[3761] <= 8'b01000000;
font_rom[3762] <= 8'b00000110;
font_rom[3763] <= 8'b01000000;
font_rom[3764] <= 8'b00000110;
font_rom[3765] <= 8'b01000000;
font_rom[3766] <= 8'b00000110;
font_rom[3767] <= 8'b01000000;
font_rom[3768] <= 8'b00000111;
font_rom[3769] <= 8'b11000000;
font_rom[3770] <= 8'b00000000;
font_rom[3771] <= 8'b00000000;
font_rom[3772] <= 8'b00000000;
font_rom[3773] <= 8'b00000000;
font_rom[3774] <= 8'b00000000;
font_rom[3775] <= 8'b00000000;
//ASCII 0x76 'v'
font_rom[3776] <= 8'b00000000;
font_rom[3777] <= 8'b00000000;
font_rom[3778] <= 8'b00000000;
font_rom[3779] <= 8'b00000000;
font_rom[3780] <= 8'b00000000;
font_rom[3781] <= 8'b00000000;
font_rom[3782] <= 8'b00000000;
font_rom[3783] <= 8'b00000000;
font_rom[3784] <= 8'b00000000;
font_rom[3785] <= 8'b00000000;
font_rom[3786] <= 8'b00000000;
font_rom[3787] <= 8'b00000000;
font_rom[3788] <= 8'b00000000;
font_rom[3789] <= 8'b00000000;
font_rom[3790] <= 8'b00000100;
font_rom[3791] <= 8'b11000000;
font_rom[3792] <= 8'b00000110;
font_rom[3793] <= 8'b11000000;
font_rom[3794] <= 8'b00000110;
font_rom[3795] <= 8'b11000000;
font_rom[3796] <= 8'b00000011;
font_rom[3797] <= 8'b10000000;
font_rom[3798] <= 8'b00000011;
font_rom[3799] <= 8'b10000000;
font_rom[3800] <= 8'b00000011;
font_rom[3801] <= 8'b00000000;
font_rom[3802] <= 8'b00000000;
font_rom[3803] <= 8'b00000000;
font_rom[3804] <= 8'b00000000;
font_rom[3805] <= 8'b00000000;
font_rom[3806] <= 8'b00000000;
font_rom[3807] <= 8'b00000000;
//ASCII 0x77 'w'
font_rom[3808] <= 8'b00000000;
font_rom[3809] <= 8'b00000000;
font_rom[3810] <= 8'b00000000;
font_rom[3811] <= 8'b00000000;
font_rom[3812] <= 8'b00000000;
font_rom[3813] <= 8'b00000000;
font_rom[3814] <= 8'b00000000;
font_rom[3815] <= 8'b00000000;
font_rom[3816] <= 8'b00000000;
font_rom[3817] <= 8'b00000000;
font_rom[3818] <= 8'b00000000;
font_rom[3819] <= 8'b00000000;
font_rom[3820] <= 8'b00000000;
font_rom[3821] <= 8'b00000000;
font_rom[3822] <= 8'b00001101;
font_rom[3823] <= 8'b11100000;
font_rom[3824] <= 8'b00001111;
font_rom[3825] <= 8'b11100000;
font_rom[3826] <= 8'b00001111;
font_rom[3827] <= 8'b11100000;
font_rom[3828] <= 8'b00001111;
font_rom[3829] <= 8'b11100000;
font_rom[3830] <= 8'b00001111;
font_rom[3831] <= 8'b11000000;
font_rom[3832] <= 8'b00000110;
font_rom[3833] <= 8'b11000000;
font_rom[3834] <= 8'b00000000;
font_rom[3835] <= 8'b00000000;
font_rom[3836] <= 8'b00000000;
font_rom[3837] <= 8'b00000000;
font_rom[3838] <= 8'b00000000;
font_rom[3839] <= 8'b00000000;
//ASCII 0x78 'x'
font_rom[3840] <= 8'b00000000;
font_rom[3841] <= 8'b00000000;
font_rom[3842] <= 8'b00000000;
font_rom[3843] <= 8'b00000000;
font_rom[3844] <= 8'b00000000;
font_rom[3845] <= 8'b00000000;
font_rom[3846] <= 8'b00000000;
font_rom[3847] <= 8'b00000000;
font_rom[3848] <= 8'b00000000;
font_rom[3849] <= 8'b00000000;
font_rom[3850] <= 8'b00000000;
font_rom[3851] <= 8'b00000000;
font_rom[3852] <= 8'b00000000;
font_rom[3853] <= 8'b00000000;
font_rom[3854] <= 8'b00001100;
font_rom[3855] <= 8'b11000000;
font_rom[3856] <= 8'b00000111;
font_rom[3857] <= 8'b11000000;
font_rom[3858] <= 8'b00000011;
font_rom[3859] <= 8'b10000000;
font_rom[3860] <= 8'b00000111;
font_rom[3861] <= 8'b00000000;
font_rom[3862] <= 8'b00001111;
font_rom[3863] <= 8'b10000000;
font_rom[3864] <= 8'b00001100;
font_rom[3865] <= 8'b11000000;
font_rom[3866] <= 8'b00000000;
font_rom[3867] <= 8'b00000000;
font_rom[3868] <= 8'b00000000;
font_rom[3869] <= 8'b00000000;
font_rom[3870] <= 8'b00000000;
font_rom[3871] <= 8'b00000000;
//ASCII 0x79 'y'
font_rom[3872] <= 8'b00000000;
font_rom[3873] <= 8'b00000000;
font_rom[3874] <= 8'b00000000;
font_rom[3875] <= 8'b00000000;
font_rom[3876] <= 8'b00000000;
font_rom[3877] <= 8'b00000000;
font_rom[3878] <= 8'b00000000;
font_rom[3879] <= 8'b00000000;
font_rom[3880] <= 8'b00000000;
font_rom[3881] <= 8'b00000000;
font_rom[3882] <= 8'b00000000;
font_rom[3883] <= 8'b00000000;
font_rom[3884] <= 8'b00000000;
font_rom[3885] <= 8'b00000000;
font_rom[3886] <= 8'b00001100;
font_rom[3887] <= 8'b01100000;
font_rom[3888] <= 8'b00001100;
font_rom[3889] <= 8'b11000000;
font_rom[3890] <= 8'b00000110;
font_rom[3891] <= 8'b11000000;
font_rom[3892] <= 8'b00000011;
font_rom[3893] <= 8'b10000000;
font_rom[3894] <= 8'b00000011;
font_rom[3895] <= 8'b10000000;
font_rom[3896] <= 8'b00000001;
font_rom[3897] <= 8'b10000000;
font_rom[3898] <= 8'b00000011;
font_rom[3899] <= 8'b00000000;
font_rom[3900] <= 8'b00000011;
font_rom[3901] <= 8'b00000000;
font_rom[3902] <= 8'b00000110;
font_rom[3903] <= 8'b00000000;
//ASCII 0x7A 'z'
font_rom[3904] <= 8'b00000000;
font_rom[3905] <= 8'b00000000;
font_rom[3906] <= 8'b00000000;
font_rom[3907] <= 8'b00000000;
font_rom[3908] <= 8'b00000000;
font_rom[3909] <= 8'b00000000;
font_rom[3910] <= 8'b00000000;
font_rom[3911] <= 8'b00000000;
font_rom[3912] <= 8'b00000000;
font_rom[3913] <= 8'b00000000;
font_rom[3914] <= 8'b00000000;
font_rom[3915] <= 8'b00000000;
font_rom[3916] <= 8'b00000000;
font_rom[3917] <= 8'b00000000;
font_rom[3918] <= 8'b00000111;
font_rom[3919] <= 8'b11100000;
font_rom[3920] <= 8'b00000000;
font_rom[3921] <= 8'b11000000;
font_rom[3922] <= 8'b00000001;
font_rom[3923] <= 8'b10000000;
font_rom[3924] <= 8'b00000001;
font_rom[3925] <= 8'b10000000;
font_rom[3926] <= 8'b00000011;
font_rom[3927] <= 8'b00000000;
font_rom[3928] <= 8'b00000111;
font_rom[3929] <= 8'b11100000;
font_rom[3930] <= 8'b00000000;
font_rom[3931] <= 8'b00000000;
font_rom[3932] <= 8'b00000000;
font_rom[3933] <= 8'b00000000;
font_rom[3934] <= 8'b00000000;
font_rom[3935] <= 8'b00000000;
//ASCII 0x7B '{'
font_rom[3936] <= 8'b00000000;
font_rom[3937] <= 8'b00000000;
font_rom[3938] <= 8'b00000000;
font_rom[3939] <= 8'b00000000;
font_rom[3940] <= 8'b00000000;
font_rom[3941] <= 8'b00000000;
font_rom[3942] <= 8'b00000000;
font_rom[3943] <= 8'b00000000;
font_rom[3944] <= 8'b00000001;
font_rom[3945] <= 8'b11000000;
font_rom[3946] <= 8'b00000011;
font_rom[3947] <= 8'b00000000;
font_rom[3948] <= 8'b00000011;
font_rom[3949] <= 8'b00000000;
font_rom[3950] <= 8'b00000011;
font_rom[3951] <= 8'b00000000;
font_rom[3952] <= 8'b00000011;
font_rom[3953] <= 8'b00000000;
font_rom[3954] <= 8'b00000111;
font_rom[3955] <= 8'b00000000;
font_rom[3956] <= 8'b00000011;
font_rom[3957] <= 8'b00000000;
font_rom[3958] <= 8'b00000011;
font_rom[3959] <= 8'b00000000;
font_rom[3960] <= 8'b00000011;
font_rom[3961] <= 8'b00000000;
font_rom[3962] <= 8'b00000011;
font_rom[3963] <= 8'b00000000;
font_rom[3964] <= 8'b00000001;
font_rom[3965] <= 8'b11000000;
font_rom[3966] <= 8'b00000000;
font_rom[3967] <= 8'b00000000;
//ASCII 0x7C '|'
font_rom[3968] <= 8'b00000000;
font_rom[3969] <= 8'b00000000;
font_rom[3970] <= 8'b00000000;
font_rom[3971] <= 8'b00000000;
font_rom[3972] <= 8'b00000000;
font_rom[3973] <= 8'b00000000;
font_rom[3974] <= 8'b00000000;
font_rom[3975] <= 8'b00000000;
font_rom[3976] <= 8'b00000001;
font_rom[3977] <= 8'b10000000;
font_rom[3978] <= 8'b00000001;
font_rom[3979] <= 8'b10000000;
font_rom[3980] <= 8'b00000001;
font_rom[3981] <= 8'b10000000;
font_rom[3982] <= 8'b00000001;
font_rom[3983] <= 8'b10000000;
font_rom[3984] <= 8'b00000001;
font_rom[3985] <= 8'b10000000;
font_rom[3986] <= 8'b00000001;
font_rom[3987] <= 8'b10000000;
font_rom[3988] <= 8'b00000001;
font_rom[3989] <= 8'b10000000;
font_rom[3990] <= 8'b00000001;
font_rom[3991] <= 8'b10000000;
font_rom[3992] <= 8'b00000001;
font_rom[3993] <= 8'b10000000;
font_rom[3994] <= 8'b00000001;
font_rom[3995] <= 8'b10000000;
font_rom[3996] <= 8'b00000001;
font_rom[3997] <= 8'b10000000;
font_rom[3998] <= 8'b00000000;
font_rom[3999] <= 8'b00000000;
//ASCII 0x7D '}'
font_rom[4000] <= 8'b00000000;
font_rom[4001] <= 8'b00000000;
font_rom[4002] <= 8'b00000000;
font_rom[4003] <= 8'b00000000;
font_rom[4004] <= 8'b00000000;
font_rom[4005] <= 8'b00000000;
font_rom[4006] <= 8'b00000000;
font_rom[4007] <= 8'b00000000;
font_rom[4008] <= 8'b00000111;
font_rom[4009] <= 8'b00000000;
font_rom[4010] <= 8'b00000001;
font_rom[4011] <= 8'b10000000;
font_rom[4012] <= 8'b00000001;
font_rom[4013] <= 8'b10000000;
font_rom[4014] <= 8'b00000001;
font_rom[4015] <= 8'b10000000;
font_rom[4016] <= 8'b00000001;
font_rom[4017] <= 8'b10000000;
font_rom[4018] <= 8'b00000001;
font_rom[4019] <= 8'b11000000;
font_rom[4020] <= 8'b00000001;
font_rom[4021] <= 8'b10000000;
font_rom[4022] <= 8'b00000001;
font_rom[4023] <= 8'b10000000;
font_rom[4024] <= 8'b00000001;
font_rom[4025] <= 8'b10000000;
font_rom[4026] <= 8'b00000001;
font_rom[4027] <= 8'b10000000;
font_rom[4028] <= 8'b00000111;
font_rom[4029] <= 8'b00000000;
font_rom[4030] <= 8'b00000000;
font_rom[4031] <= 8'b00000000;
//ASCII 0x7E '~'
font_rom[4032] <= 8'b00000000;
font_rom[4033] <= 8'b00000000;
font_rom[4034] <= 8'b00000000;
font_rom[4035] <= 8'b00000000;
font_rom[4036] <= 8'b00000000;
font_rom[4037] <= 8'b00000000;
font_rom[4038] <= 8'b00000000;
font_rom[4039] <= 8'b00000000;
font_rom[4040] <= 8'b00000000;
font_rom[4041] <= 8'b00000000;
font_rom[4042] <= 8'b00000000;
font_rom[4043] <= 8'b00000000;
font_rom[4044] <= 8'b00000000;
font_rom[4045] <= 8'b00000000;
font_rom[4046] <= 8'b00000111;
font_rom[4047] <= 8'b01000000;
font_rom[4048] <= 8'b00001111;
font_rom[4049] <= 8'b11000000;
font_rom[4050] <= 8'b00001101;
font_rom[4051] <= 8'b11000000;
font_rom[4052] <= 8'b00000000;
font_rom[4053] <= 8'b00000000;
font_rom[4054] <= 8'b00000000;
font_rom[4055] <= 8'b00000000;
font_rom[4056] <= 8'b00000000;
font_rom[4057] <= 8'b00000000;
font_rom[4058] <= 8'b00000000;
font_rom[4059] <= 8'b00000000;
font_rom[4060] <= 8'b00000000;
font_rom[4061] <= 8'b00000000;
font_rom[4062] <= 8'b00000000;
font_rom[4063] <= 8'b00000000;
//ASCII 0x7F ''
font_rom[4064] <= 8'b00000000;
font_rom[4065] <= 8'b00000000;
font_rom[4066] <= 8'b00000000;
font_rom[4067] <= 8'b00000000;
font_rom[4068] <= 8'b00000000;
font_rom[4069] <= 8'b00000000;
font_rom[4070] <= 8'b00000000;
font_rom[4071] <= 8'b00000000;
font_rom[4072] <= 8'b00000011;
font_rom[4073] <= 8'b10000000;
font_rom[4074] <= 8'b00000010;
font_rom[4075] <= 8'b10000000;
font_rom[4076] <= 8'b00000010;
font_rom[4077] <= 8'b10000000;
font_rom[4078] <= 8'b00000010;
font_rom[4079] <= 8'b10000000;
font_rom[4080] <= 8'b00000010;
font_rom[4081] <= 8'b10000000;
font_rom[4082] <= 8'b00000010;
font_rom[4083] <= 8'b10000000;
font_rom[4084] <= 8'b00000010;
font_rom[4085] <= 8'b10000000;
font_rom[4086] <= 8'b00000011;
font_rom[4087] <= 8'b10000000;
font_rom[4088] <= 8'b00000000;
font_rom[4089] <= 8'b00000000;
font_rom[4090] <= 8'b00000000;
font_rom[4091] <= 8'b00000000;
font_rom[4092] <= 8'b00000000;
font_rom[4093] <= 8'b00000000;
font_rom[4094] <= 8'b00000000;
font_rom[4095] <= 8'b00000000;


always @(posedge clk) begin
	out <= font_rom[address];
end

endmodule