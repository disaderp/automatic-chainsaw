module Buff(
	input clk,
	